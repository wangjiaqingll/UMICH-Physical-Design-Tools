LAYER met1
     TYPE ROUTING ;
     WIDTH 0.2 ;
     OFFSET 0.00 ;
     PITCH 0.7 ;
     SPACING 0.2 RANGE 0.1 10.0 ;
     SPACING 0.60 RANGE 10 35 ;
     DIRECTION HORIZONTAL ;
     CAPACITANCE CPERSQDIST 5.0e-05 ;
     EDGECAPACITANCE 6.0e-05 ;
     RESISTANCE RPERSQ 0.1 ;
     CAPMULTIPLIER 1.00 ;
END met1

