#CREATE TIME 31 March 1994 15:30:41
NAMESCASESENSITIVE OFF ;
#TECHNOLOGY SECTION

LAYER PWELL
  TYPE MASTERSLICE ;
END PWELL

LAYER NDIFF
  TYPE MASTERSLICE ;
END NDIFF

LAYER PDIFF
  TYPE MASTERSLICE ;
END PDIFF

LAYER POLY
  TYPE MASTERSLICE ;
END POLY

LAYER CONT
  TYPE CUT ;
END CONT

LAYER MET1
  TYPE ROUTING ;
  PITCH 4.8 ;
  WIDTH 1.6 ;
  SPACING 1.4 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ .8E-01 ;
  CAPACITANCE CPERSQDIST .192E-03 ;
END MET1

LAYER VIA
  TYPE CUT ;
END VIA

LAYER MET2
  TYPE ROUTING ;
  PITCH 4.8 ;
  WIDTH 2 ;
  SPACING 1.6 ;
  DIRECTION VERTICAL ;
  RESISTANCE RPERSQ .32E-01 ;
  CAPACITANCE CPERSQDIST .88E-04 ;
END MET2

VIA M1M2 DEFAULT 
  LAYER MET1 ;
    RECT -1.7 -1.7 1.7 1.7 ;
  LAYER VIA ;
    RECT -.7 -.7 .7 .7 ;
  LAYER MET2 ;
    RECT -1.6 -1.6 1.6 1.6 ;
END M1M2
VIA PMET1 DEFAULT 
  LAYER POLY ;
    RECT -1.4 -1.4 1.4 1.4 ;
  LAYER CONT ;
    RECT -.6 -.6 .6 .6 ;
  LAYER MET1 ;
    RECT -1.4 -1.4 1.4 1.4 ;
END PMET1
VIA BIGM1M2
  LAYER MET1 ;
    RECT -1.7 -1.7 1.7 1.7 ;
  LAYER VIA ;
    RECT -.7 -.7 .7 .7 ;
  LAYER MET2 ;
    RECT -1.6 -1.6 1.6 1.6 ;
END BIGM1M2

SPACING
  SAMENET VIA POLY 1 ;
  SAMENET CONT CONT 1.4 ;
  SAMENET VIA CONT 1.6 ;
  SAMENET VIA VIA 1 ;
END SPACING

#SITE SECTION
SITE CORE
  SIZE 4.8 BY 36.8 ;
  CLASS CORE ;
END CORE

SITE CORE1
  SIZE 958.1 BY 150 ;
  CLASS CORE ;
END CORE1

SITE IO
  SIZE 3.6 BY 3.6 ;
  CLASS PAD ;
END IO

#MACRO SECTION

MACRO DUMMY_1 
  CLASS CORE ;
  SIZE 9.6 BY 36.8 ;
  ORIGIN 0 0 ;
  SYMMETRY X  ;
  SITE CORE 0 0 N DO 1 BY 1 STEP 0 0 ;
  PIN O
  DIRECTION OUTPUT ;
  USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT .8 9.3 4.1 22.7 ;
    END
  END O
  PIN I
  DIRECTION INPUT ;
  USE SIGNAL ;
  CAPACITANCE .3312E-01 ;
    PORT
      LAYER POLY ;
        RECT .6 -5 4.2 -1.4 ;
    END
    PORT
      LAYER POLY ;
        RECT 5.4 14.2 9 17.8 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 43 4.2 46.6 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 47.8 4.2 51.4 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 -14.6 4.2 -11 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 38.2 4.2 41.8 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 -9.8 4.2 -6.2 ;
    END
  END I
  PIN VSS
  DIRECTION INOUT ;
  SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.6 3.2 ;
    END
  END VSS
  PIN VCC
  DIRECTION INOUT ;
  SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 33.6 9.6 36.8 ;
    END
  END VCC
  OBS
      LAYER VIA ;
      RECT 4.3 14.1 5.4 17.9 ;
      RECT 4.3 17.9 5.3 34.5 ;
      RECT 4.3 5.1 5.3 14.1 ;
      RECT 6.6 1 7.8 2.2 ;
      RECT 6.6 34.6 7.8 35.8 ;
      RECT 2.1 10.1 3.3 11.3 ;
      RECT 2.1 20.7 3.3 21.9 ;
  END
  TIMING
   FROMPIN  I  ;    TOPIN  O  ;  
    RISE INTRINSIC  .109 .109 VARIABLE 2.1957 2.1957 ;
    FALL INTRINSIC  .121 .121 VARIABLE 2.432 2.432 ;
    UNATENESS INVERT ;
  END TIMING
END DUMMY_1 

MACRO DUMMY_2 
  CLASS CORE ;
  SIZE 14.4 BY 36.8 ;
  ORIGIN 0 0 ;
  SYMMETRY X  ;
  SITE CORE 0 0 N DO 1 BY 1 STEP 0 0 ;
  PIN O
  DIRECTION OUTPUT ;
  USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT .8 9.3 5.6 12.8 ;
        RECT 5.6 9.3 8.8 22.7 ;
    END
  END O
  PIN I2
  DIRECTION INPUT ;
  USE SIGNAL ;
  CAPACITANCE .2208E-01 ;
    PORT
      LAYER POLY ;
        RECT 10.2 38.2 13.8 41.8 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 -9.8 13.8 -6.2 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 14.2 13.8 17.8 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 -5 13.8 -1.4 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 43 13.8 46.6 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 47.8 13.8 51.4 ;
    END
    PORT
      LAYER POLY ;
        RECT 10.2 -14.6 13.8 -11 ;
    END
  END I2
  PIN I1
  DIRECTION INPUT ;
  USE SIGNAL ;
  CAPACITANCE .2208E-01 ;
    PORT
      LAYER POLY ;
        RECT .6 -5 4.2 -1.4 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 47.8 4.2 51.4 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 38.2 4.2 41.8 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 43 4.2 46.6 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 -14.6 4.2 -11 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 -9.8 4.2 -6.2 ;
    END
    PORT
      LAYER POLY ;
        RECT .6 14.2 4.2 17.8 ;
    END
  END I1
  PIN VSS
  DIRECTION INOUT ;
  SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.4 3.2 ;
    END
  END VSS
  PIN VCC
  DIRECTION INOUT ;
  SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 33.6 14.4 36.8 ;
    END
  END VCC
  OBS
      LAYER VIA ;
      RECT 9.1 14.1 10.2 17.9 ;
      RECT 9.1 17.9 10.1 27.5 ;
      RECT 9.1 5.1 10.1 14.1 ;
      RECT 4.3 17.9 5.3 27.5 ;
      RECT 4.3 5.1 5.3 14.1 ;
      RECT 4.2 14.1 5.3 17.9 ;
      RECT 11.4 1 12.6 2.2 ;
      RECT 11.4 34.6 12.6 35.8 ;
      RECT 1.8 34.6 3 35.8 ;
      RECT 6.6 20.7 7.8 21.9 ;
      RECT 2.1 10.1 3.3 11.3 ;
  END
  TIMING
   FROMPIN  I1  I2  ;    TOPIN  O  ;  
    RISE INTRINSIC  .293 .293 VARIABLE 4.7424 4.7424 ;
    FALL INTRINSIC  .127 .127 VARIABLE 3.8037 3.8037 ;
    UNATENESS INVERT ;
  END TIMING
END DUMMY_2

MACRO IOCELL
  CLASS PAD ;
  SIZE 3.6 BY 3.6 ;
  ORIGIN 0 0 ;
  SYMMETRY R90  ;
  SITE IO 0 0 N DO 1 BY 1 STEP 0 0 ;
  PIN IN
  DIRECTION INOUT ;
  USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT .8 .8 2.8 2.8 ;
    END
  END IN
END IOCELL

MACRO IOCELL1
  CLASS PAD ;
  SIZE 3.6 BY 3.6 ;
  ORIGIN 0 0 ;
  SYMMETRY R90  ;
  SITE IO 0 0 N DO 1 BY 1 STEP 0 0 ;
  PIN IN
  DIRECTION INOUT ;
  USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT .8 .8 2.8 2.8 ;
    END
  END IN
END IOCELL1

END LIBRARY
