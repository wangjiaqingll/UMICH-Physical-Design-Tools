#
# CMOS26G LEF technology file
# @(#) 1.3 92/08/12  13:40:42   Eric A. Slutz
#
#       Updated         05/12/93    sjr
#       Updated         06/08/93    sjr
#       Updated         06/09/93    sjr
#       Updated         07/07/93    sjr
#       Modified manually to add the old 26R pads and site types - by
#       Modifed manually to add the corrected TRIZDD cell (08/06/83) - by
#       Modified manually to add case sensitive names (8/17/93) - by
# 
#############################################################################

NAMESCASESENSITIVE ON ;

#Note: no other values are allowed at this time
#  all commented out so that a warning is not generated.
#UNITS
  # not allowed in lef: DISTANCE MICRON 1 ;
#  TIME NANOSECONDS 1 ;
#  CAPACITANCE PICOFARADS 1 ;
#  RESISTANCE OHMS 1 ;
#  POWER MILLIWATTS 1 ;
#  CURRENT MILLIAMPS 1 ;
#  VOLTAGE VOLTS 1 ;
#END UNITS

LAYER poly
# no routing will be done in poly
  TYPE MASTERSLICE ;
END poly

LAYER cont1
  TYPE CUT ;
END cont1

LAYER metal1
  TYPE ROUTING ; PITCH 2.4 ; WIDTH 1.0 ; SPACING 1.0 ;
  DIRECTION HORIZONTAL ; 
# timing analysis
  RESISTANCE RPERSQ .090 ; # max at 85C
# CAPACITANCE CPERSQDIST .000235 ; # per square micron (max)
  CAPACITANCE CPERSQDIST .000195 ; # per square micron (nom)
#                                   Hive generated, M1 arrays above sub under
#                                   M2. w=1.0um sp=1.2um & M1 arrays above
#                                   poly under M2. w=1.0um sp=1.2um.
# more accurate model
  #eas HEIGHT 0.0 ;
  #eas THICKNESS 0.0 ;
  #eas SHRINKAGE 0.0 ;
  #eas CAPMULTIPLIER 1.0 ;
END metal1

LAYER cont2
  TYPE CUT ; 
END cont2

LAYER metal2
  TYPE ROUTING ; PITCH 2.6 ; WIDTH 1.0 ; SPACING 1.0 ;
  DIRECTION VERTICAL ;
# timing analysis
  RESISTANCE RPERSQ .090 ; # max at 85C
# CAPACITANCE CPERSQDIST .000235 ; # per square micron (max)
  CAPACITANCE CPERSQDIST .000185 ; # per square micron (nom)
#                                    Hive generated, M2 arrays above sub, under
#                                    M3 plane. w=1.0um, sp=1.2um & M2 arrays
#                                    above sparse M1 & sub, under M3
#                                    w=1.0um, sp=1.2um.
END metal2

LAYER cont3
  TYPE CUT ;
END cont3

LAYER metal3
  TYPE ROUTING ; PITCH 3.2 ; WIDTH 1.8 ; SPACING 1.2 ;
  DIRECTION HORIZONTAL ;
# timing analysis
  RESISTANCE RPERSQ .065 ; # max at 85C
# CAPACITANCE CPERSQDIST .000120 ; # per square micron (max)
  CAPACITANCE CPERSQDIST .000100 ; # per square micron (nom)
#                                    Hive generated, M3 arrays above M2 + M1
#                                    plane-averaged. w=1.8um, sp=1.7um
END metal3

VIA via01 DEFAULT
  #eas FOREIGN VIA01 0 0 ;
  LAYER poly      ; RECT -0.8 -0.8 0.8 0.8 ; # 8A1 & 8G
  LAYER cont1     ; RECT -0.4 -0.4 0.4 0.4 ; # 8A1
  LAYER metal1    ; RECT -0.8 -0.8 0.8 0.8 ; # 8A1 & 8E1
  RESISTANCE 8.0 ; # nom at 110C
END via01

VIA via12 DEFAULT
  LAYER metal1    ; RECT -0.8 -0.8 0.8 0.8 ; # 10A1 & 10D
  LAYER cont2     ; RECT -0.4 -0.4 0.4 0.4 ; # 10A1 
  LAYER metal2    ; RECT -0.8 -0.8 0.8 0.8 ; # 10A1 & 10E
  RESISTANCE 1.5 ; # max at 110C
END via12

VIA via23 DEFAULT
  LAYER metal2    ; RECT -0.8 -0.8 0.8 0.8 ; # 12A1 & 12D
  LAYER cont3     ; RECT -0.4 -0.4 0.4 0.4 ; # 12A1
  LAYER metal3    ; RECT -1.0 -1.0 1.0 1.0 ; # 12A1 & 12E
  RESISTANCE 1.5 ; # max at 110C
END via23

VIA stripevia
  FOREIGN ZZSTRVIA68 ;
  layer metal1   ; rect -3.4 -2.8  3.4 2.8 ;
  layer metal2   ; rect -3.4 -2.8  3.4 2.8 ;
  layer cont2    ; rect -2.4 -0.4 -1.6 0.4 ;
                   rect -0.4 -0.4  0.4 0.4 ;
                   rect  1.6 -0.4  2.4 0.4 ;
END stripevia

VIARULE turnm1 GENERATE
   LAYER metal1 ; DIRECTION VERTICAL ;
   LAYER metal1 ; DIRECTION HORIZONTAL ;
END turnm1

VIARULE turnm2 GENERATE
   LAYER metal2 ; DIRECTION VERTICAL ;
   LAYER metal2 ; DIRECTION HORIZONTAL ;
END turnm2

VIARULE turnm3 GENERATE
   LAYER metal3 ; DIRECTION VERTICAL ;
   LAYER metal3 ; DIRECTION HORIZONTAL ;
END turnm3

VIARULE pwrstripe
  layer metal1 ; direction horizontal ; width 5.6 to 5.6 ;
  layer metal2 ; direction vertical ; width 6.8 to 6.8 ;
  via stripevia ;
END pwrstripe

VIARULE array12 GENERATE
  LAYER metal1 ; DIRECTION horizontal ;
    OVERHANG 0.4 ; # Rule 10D
  LAYER metal2 ; DIRECTION vertical ;
    OVERHANG 0.4 ; # Rule 10E
  LAYER cont2 ;
    RECT -0.4 -0.4 0.4 0.4 ; # Rule 10A1
    SPACING 2.0 BY 2.0 ; # Rule 10A1 & 10B
  RESISTANCE 1.5 ;
END array12

VIARULE array23 GENERATE
  LAYER metal2 ; DIRECTION vertical ;
    OVERHANG 0.6 ; # Rule 12D  (modified to get around a Cell problem - by)
  LAYER metal3 ; DIRECTION horizontal ;
    OVERHANG 0.6 ; # Rule 12E
  LAYER cont3 ;
    RECT -0.4 -0.4 0.4 0.4 ; # Rule 12A
    SPACING 2.0 BY 2.0 ; # Rule 12A1 & 12B
  RESISTANCE 1.5 ;
END array23

SPACING
  SAMENET cont2 cont2 1.2 ; # Rule 10B
  SAMENET cont1 cont2 0.6 ; # Rule 10C1
  SAMENET cont3 cont3 1.2 ; # Rule 12B
  SAMENET cont2 cont3 0.6 ; # Rule 12C
END SPACING

#eas IRDROP

#eas MINFEATURE

#eas DIELECTRIC

SITE CORE26  CLASS CORE ; SYMMETRY    Y ; SIZE   2.6 BY  38.4 ; END CORE26
#Site for dummy IO ports
SITE SMALLIO  CLASS PAD ;                SIZE   1.3 BY   1.3 ; END SMALLIO

# Pad site.  Need to have 5.2um wide site to allow even insertion of
# ZZPADSPC cells
site target      CLASS PAD ; size   5.2 by 551.2 ;          end target

# Corner sites
site nwcorner    CLASS PAD ; size 551.2 by 551.2 ;    end nwcorner
site necorner    CLASS PAD ; size 551.2 by 551.2 ;    end necorner
site secorner    CLASS PAD ; size 551.2 by 551.2 ;  end secorner
site swcorner    CLASS PAD ; size 551.2 by 551.2 ;  end swcorner

MACRO AND2EE
  CLASS CORE ;
  FOREIGN AND2EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 3.400 6.700 4.400 17.300 ;
      RECT 3.400 16.300 7.000 17.300 ;
      RECT 6.000 16.300 7.000 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 3.400 11.500 9.600 12.500 ;
      RECT 3.400 16.300 7.000 19.700 ;
      RECT 0.800 18.700 7.000 19.700 ;
      RECT 3.400 23.500 9.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
  END
END AND2EE

MACRO AND2FF
  CLASS CORE ;
  FOREIGN AND2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 10.100 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 18.700 7.000 19.700 ;
      RECT 6.000 18.700 7.000 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 3.400 6.700 4.400 24.500 ;
      RECT 3.400 11.500 9.600 12.500 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 3.400 18.700 7.000 22.100 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
  END
END AND2FF

MACRO AND2GG
  CLASS CORE ;
  FOREIGN AND2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 17.300 ; # Q|0.0@0
      RECT 0.800 16.300 4.400 17.300 ; # Q|0.0@1
      RECT 3.400 16.300 4.400 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 3.400 6.700 4.400 14.900 ;
      RECT 3.400 13.900 9.600 14.900 ;
      RECT 8.600 13.900 9.600 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 0.800 4.300 12.200 7.700 ;
      RECT 0.800 4.300 7.000 10.100 ;
      RECT 3.400 4.300 4.400 19.700 ;
      RECT 11.200 11.500 12.200 12.500 ;
      RECT 3.400 13.900 9.600 14.900 ;
      RECT 8.600 13.900 9.600 19.700 ;
      RECT 0.800 18.700 4.400 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END AND2GG

MACRO AND2HH
  CLASS CORE ;
  FOREIGN AND2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 6.000 18.700 9.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 3.400 4.300 12.200 7.700 ;
      RECT 3.400 4.300 9.600 10.100 ;
      RECT 6.000 11.500 12.200 12.500 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 3.400 16.300 9.600 19.700 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END AND2HH

MACRO AND3EE
  CLASS CORE ;
  FOREIGN AND3EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 6.000 18.700 9.600 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 12.200 5.300 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 12.200 7.700 ;
      RECT 6.000 4.300 7.000 22.100 ;
      RECT 11.200 4.300 12.200 10.100 ;
      RECT 3.400 11.500 7.000 17.300 ;
      RECT 3.400 13.900 12.200 17.300 ;
      RECT 0.800 16.300 12.200 17.300 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 13.900 9.600 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 13.900 9.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
  END
END AND3EE

MACRO AND3FF
  CLASS CORE ;
  FOREIGN AND3FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 6.000 18.700 9.600 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 12.200 5.300 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 12.200 7.700 ;
      RECT 6.000 4.300 7.000 22.100 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 6.000 13.900 12.200 17.300 ;
      RECT 0.800 18.700 1.800 19.700 ;
      RECT 6.000 13.900 9.600 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 23.500 12.200 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 12.200 29.300 ;
  END
END AND3FF

MACRO AND3GG
  CLASS CORE ;
  FOREIGN AND3GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 16.300 12.200 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 7.700 ; # Q|0.0@0
      RECT 0.800 9.100 1.800 17.300 ; # Q|0.0@1
      RECT 3.400 18.700 4.400 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 9.100 7.000 17.300 ;
      RECT 11.200 11.500 12.200 14.900 ;
      RECT 3.400 16.300 9.600 17.300 ;
      RECT 6.000 18.700 14.800 19.700 ;
      RECT 13.800 18.700 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 13.800 4.300 14.800 5.300 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 11.200 11.500 12.200 14.900 ;
      RECT 11.200 13.900 14.800 14.900 ;
      RECT 0.800 16.300 9.600 19.700 ;
      RECT 13.800 13.900 14.800 22.100 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 12.200 29.300 ;
  END
END AND3GG

MACRO AND3HH
  CLASS CORE ;
  FOREIGN AND3HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 10.100 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 14.900 ; # Q|0.0@0
      RECT 3.400 18.700 4.400 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 14.800 7.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 6.000 11.500 9.600 17.300 ;
      RECT 6.000 13.900 12.200 17.300 ;
      RECT 0.800 16.300 12.200 17.300 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 8.600 18.700 14.800 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 7.000 5.300 ;
      RECT 13.800 4.300 14.800 10.100 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 8.600 6.700 14.800 7.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 6.000 11.500 9.600 17.300 ;
      RECT 6.000 13.900 14.800 17.300 ;
      RECT 0.800 16.300 14.800 17.300 ;
      RECT 0.800 16.300 4.400 19.700 ;
      RECT 8.600 13.900 14.800 19.700 ;
      RECT 13.800 13.900 14.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END AND3HH

MACRO AND4EE
  CLASS CORE ;
  FOREIGN AND4EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 14.800 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 6.000 16.300 14.800 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 13.800 4.300 14.800 7.700 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 6.700 14.800 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 13.900 14.800 14.900 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 13.900 14.800 19.700 ;
      RECT 3.400 23.500 9.600 24.500 ;
  END
END AND4EE

MACRO AND4FF
  CLASS CORE ;
  FOREIGN AND4FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 14.800 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 6.000 18.700 14.800 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 14.800 7.700 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 6.000 16.300 14.800 19.700 ;
      RECT 0.800 18.700 1.800 19.700 ;
      RECT 11.200 16.300 14.800 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
  END
END AND4FF

MACRO AND4GG
  CLASS CORE ;
  FOREIGN AND4GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 10.100 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 14.800 7.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 12.200 10.100 ;
      RECT 3.400 11.500 7.000 17.300 ;
      RECT 3.400 13.900 12.200 17.300 ;
      RECT 0.800 18.700 4.400 19.700 ;
      RECT 8.600 13.900 12.200 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 0.800 4.300 4.400 10.100 ;
      RECT 11.200 4.300 14.800 10.100 ;
      RECT 0.800 6.700 14.800 7.700 ;
      RECT 8.600 6.700 14.800 10.100 ;
      RECT 3.400 11.500 7.000 17.300 ;
      RECT 3.400 13.900 12.200 17.300 ;
      RECT 0.800 18.700 4.400 19.700 ;
      RECT 8.600 13.900 12.200 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 14.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 14.800 29.300 ;
  END
END AND4GG

MACRO AND4HH
  CLASS CORE ;
  FOREIGN AND4HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 13.900 17.400 17.300 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 17.300 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 17.300 ; # Q|0.0@0
      RECT 3.400 18.700 4.400 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 6.000 18.700 14.800 22.100 ;
      RECT 3.400 21.100 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 7.000 7.700 ;
      RECT 16.400 4.300 17.400 10.100 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 3.400 4.300 7.000 22.100 ;
      RECT 3.400 11.500 9.600 12.500 ;
      RECT 11.200 13.900 17.400 14.900 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 3.400 18.700 14.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 18.700 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END AND4HH

MACRO AOI211DD
  CLASS CORE ;
  FOREIGN AOI211DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 7.700 ; # Q|0.0@0
      RECT 21.600 6.700 22.600 17.300 ; # Q|0.0@1
      RECT 3.400 16.300 4.400 17.300 ; # Q|0.0@2
      RECT 8.600 16.300 9.600 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 20.000 10.100 ;
      RECT 6.000 9.100 20.000 10.100 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 8.600 6.700 14.800 12.500 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 19.000 13.900 20.000 19.700 ;
      RECT 6.000 16.300 7.000 19.700 ;
      RECT 11.200 16.300 20.000 19.700 ;
      RECT 0.800 18.700 22.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 22.600 5.300 ;
      RECT 3.400 6.700 20.000 7.700 ;
      RECT 6.000 4.300 20.000 10.100 ;
      RECT 0.800 11.500 4.400 12.500 ;
      RECT 8.600 4.300 20.000 12.500 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 16.400 4.300 20.000 19.700 ;
      RECT 0.800 16.300 7.000 19.700 ;
      RECT 11.200 16.300 22.600 19.700 ;
      RECT 0.800 18.700 22.600 19.700 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 6.000 13.900 7.000 22.100 ;
      RECT 16.400 4.300 17.400 22.100 ;
      RECT 21.600 16.300 22.600 22.100 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END AOI211DD

MACRO AOI211FF
  CLASS CORE ;
  FOREIGN AOI211FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 33.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
      RECT 11.200 9.100 14.800 10.100 ; # A|0.0@1
      RECT 21.600 9.100 22.600 10.100 ; # A|0.0@2
      RECT 29.400 9.100 30.400 10.100 ; # A|0.0@3
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 13.900 25.200 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 6.700 33.000 17.300 ; # Q|0.0@0
      RECT 3.400 16.300 14.800 17.300 ; # Q|0.0@1
      RECT 26.800 16.300 27.800 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 33.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 33.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 30.400 7.700 ;
      RECT 6.000 6.700 9.600 10.100 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 24.200 6.700 27.800 12.500 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 8.600 11.500 30.400 12.500 ;
      RECT 11.200 11.500 22.600 14.900 ;
      RECT 29.400 11.500 30.400 22.100 ;
      RECT 16.400 16.300 25.200 22.100 ;
      RECT 0.800 18.700 33.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 24.200 -0.500 27.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 33.000 5.300 ;
      RECT 6.000 4.300 30.400 7.700 ;
      RECT 6.000 4.300 9.600 10.100 ;
      RECT 16.400 4.300 20.000 22.100 ;
      RECT 24.200 4.300 27.800 12.500 ;
      RECT 0.800 11.500 4.400 22.100 ;
      RECT 8.600 11.500 30.400 12.500 ;
      RECT 0.800 13.900 22.600 14.900 ;
      RECT 29.400 11.500 30.400 22.100 ;
      RECT 16.400 16.300 25.200 22.100 ;
      RECT 0.800 18.700 33.000 22.100 ;
      RECT 11.200 18.700 12.200 24.500 ;
      RECT 21.600 11.500 22.600 24.500 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END AOI211FF

MACRO AOI21DD
  CLASS CORE ;
  FOREIGN AOI21DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 3.400 6.700 4.400 12.500 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 18.700 9.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 8.600 4.300 9.600 5.300 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 3.400 6.700 4.400 12.500 ;
      RECT 8.600 11.500 9.600 12.500 ;
      RECT 0.800 13.900 1.800 14.900 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 0.800 18.700 9.600 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END AOI21DD

MACRO AOI21FF
  CLASS CORE ;
  FOREIGN AOI21FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 4.400 10.100 ; # C|0.0@0
      RECT 11.200 9.100 12.200 10.100 ; # C|0.0@1
      RECT 13.800 11.500 14.800 12.500 ; # C|0.0@2
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 6.700 12.200 7.700 ; # Q|0.0@0
      RECT 16.400 6.700 17.400 17.300 ; # Q|0.0@1
      RECT 6.000 16.300 7.000 17.300 ; # Q|0.0@2
      RECT 11.200 16.300 12.200 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 7.700 ;
      RECT 6.000 6.700 9.600 10.100 ;
      RECT 13.800 6.700 14.800 10.100 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 13.800 16.300 14.800 22.100 ;
      RECT 3.400 18.700 17.400 19.700 ;
      RECT 3.400 18.700 14.800 22.100 ;
    LAYER cont2 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 6.000 4.300 17.400 5.300 ;
      RECT 6.000 4.300 9.600 12.500 ;
      RECT 13.800 4.300 17.400 7.700 ;
      RECT 0.800 9.100 9.600 10.100 ;
      RECT 13.800 4.300 14.800 10.100 ;
      RECT 3.400 16.300 14.800 22.100 ;
      RECT 0.800 18.700 17.400 19.700 ;
      RECT 0.800 18.700 14.800 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END AOI21FF

MACRO AOI221DD
  CLASS CORE ;
  FOREIGN AOI221DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 25.200 10.100 ; # A|0.0@0
      RECT 13.800 9.100 14.800 12.500 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 11.500 27.800 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 10.100 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 11.500 30.400 14.900 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 17.300 ; # Q|0.0@0
      RECT 11.200 6.700 20.000 7.700 ; # Q|0.0@1
      RECT 6.000 16.300 9.600 17.300 ; # Q|0.0@2
      RECT 24.200 16.300 25.200 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 7.700 ;
      RECT 21.600 6.700 25.200 7.700 ;
      RECT 8.600 11.500 12.200 12.500 ;
      RECT 24.200 11.500 25.200 14.900 ;
      RECT 11.200 16.300 22.600 22.100 ;
      RECT 29.400 16.300 30.400 19.700 ;
      RECT 0.800 18.700 30.400 19.700 ;
      RECT 8.600 18.700 27.800 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 16.400 -0.500 20.000 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 3.400 4.300 25.200 5.300 ;
      RECT 29.400 4.300 30.400 5.300 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 21.600 4.300 25.200 7.700 ;
      RECT 11.200 9.100 12.200 24.500 ;
      RECT 24.200 4.300 25.200 24.500 ;
      RECT 3.400 11.500 4.400 12.500 ;
      RECT 8.600 11.500 12.200 14.900 ;
      RECT 16.400 11.500 25.200 24.500 ;
      RECT 8.600 13.900 25.200 14.900 ;
      RECT 29.400 13.900 30.400 19.700 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 6.000 16.300 7.000 22.100 ;
      RECT 11.200 13.900 25.200 24.500 ;
      RECT 0.800 18.700 30.400 19.700 ;
      RECT 6.000 18.700 27.800 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 18.700 27.800 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
  END
END AOI221DD

MACRO AOI222DD
  CLASS CORE ;
  FOREIGN AOI222DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 39.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 11.500 30.400 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 11.500 33.000 14.900 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # E|0.0@0
    END
  END E
  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 22.600 10.100 ; # F|0.0@0
      RECT 29.400 9.100 35.600 10.100 ; # F|0.0@1
      RECT 34.600 9.100 35.600 14.900 ; # F|0.0@2
    END
  END F
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 17.400 7.700 ; # Q|0.0@1
      RECT 3.400 6.700 4.400 17.300 ; # Q|0.0@2
      RECT 3.400 16.300 7.000 17.300 ; # Q|0.0@3
      RECT 13.800 16.300 27.800 17.300 ; # Q|0.0@4
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 39.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 39.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 11.200 6.700 12.200 7.700 ;
      RECT 19.000 6.700 27.800 7.700 ;
      RECT 24.200 6.700 27.800 12.500 ;
      RECT 19.000 11.500 27.800 12.500 ;
      RECT 8.600 13.900 22.600 14.900 ;
      RECT 8.600 13.900 12.200 22.100 ;
      RECT 3.400 18.700 35.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 0.800 4.300 27.800 5.300 ;
      RECT 32.000 4.300 33.000 7.700 ;
      RECT 6.000 4.300 7.000 7.700 ;
      RECT 11.200 4.300 12.200 24.500 ;
      RECT 19.000 6.700 35.600 7.700 ;
      RECT 24.200 4.300 27.800 14.900 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 11.200 11.500 27.800 14.900 ;
      RECT 34.600 11.500 35.600 12.500 ;
      RECT 8.600 13.900 33.000 14.900 ;
      RECT 8.600 13.900 12.200 24.500 ;
      RECT 26.800 13.900 30.400 24.500 ;
      RECT 0.800 18.700 35.600 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 6.000 18.700 33.000 24.500 ;
      RECT 37.200 23.500 38.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
  END
END AOI222DD

MACRO AOI222FF
  CLASS CORE ;
  FOREIGN AOI222FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 57.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 9.100 53.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 45.000 9.100 46.000 14.900 ; # B|0.0@0
      RECT 32.000 13.900 35.600 14.900 ; # B|0.0@1
      RECT 42.400 13.900 46.000 14.900 ; # B|0.0@2
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 9.100 40.800 12.500 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # E|0.0@0
    END
  END E
  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 10.100 ; # F|0.0@0
      RECT 37.200 9.100 38.200 10.100 ; # F|0.0@1
    END
  END F
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 14.800 7.700 ; # Q|0.0@1
      RECT 42.400 6.700 56.400 7.700 ; # Q|0.0@2
      RECT 55.400 6.700 56.400 17.300 ; # Q|0.0@3
      RECT 29.400 16.300 43.400 17.300 ; # Q|0.0@4
      RECT 47.600 16.300 56.400 17.300 ; # Q|0.0@5
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 57.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 57.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 12.200 22.100 ;
      RECT 16.400 6.700 40.800 7.700 ;
      RECT 16.400 6.700 35.600 12.500 ;
      RECT 3.400 11.500 38.200 12.500 ;
      RECT 0.800 13.900 30.400 14.900 ;
      RECT 37.200 13.900 40.800 14.900 ;
      RECT 8.600 11.500 27.800 22.100 ;
      RECT 45.000 16.300 46.000 22.100 ;
      RECT 3.400 18.700 53.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 32.000 -0.500 35.600 0.500 ;
      RECT 47.600 -0.500 51.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 56.400 5.300 ;
      RECT 6.000 4.300 12.200 7.700 ;
      RECT 16.400 4.300 43.400 7.700 ;
      RECT 8.600 4.300 12.200 24.500 ;
      RECT 16.400 4.300 35.600 12.500 ;
      RECT 52.800 9.100 53.800 10.100 ;
      RECT 0.800 11.500 40.800 12.500 ;
      RECT 45.000 11.500 46.000 12.500 ;
      RECT 0.800 11.500 30.400 14.900 ;
      RECT 37.200 11.500 40.800 14.900 ;
      RECT 8.600 11.500 27.800 24.500 ;
      RECT 45.000 16.300 48.600 24.500 ;
      RECT 0.800 18.700 56.400 19.700 ;
      RECT 0.800 18.700 53.800 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 6.000 18.700 48.600 24.500 ;
      RECT 55.400 23.500 56.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 55.400 28.300 56.400 29.300 ;
  END
END AOI222FF

MACRO AOI22DD
  CLASS CORE ;
  FOREIGN AOI22DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 12.500 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 17.300 ; # Q|0.0@0
      RECT 6.000 16.300 9.600 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 3.400 6.700 4.400 12.500 ;
      RECT 6.000 13.900 7.000 14.900 ;
      RECT 3.400 18.700 9.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 6.000 4.300 9.600 5.300 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 0.800 6.700 4.400 12.500 ;
      RECT 11.200 11.500 12.200 12.500 ;
      RECT 6.000 13.900 7.000 22.100 ;
      RECT 0.800 18.700 9.600 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END AOI22DD

MACRO AOI22FF
  CLASS CORE ;
  FOREIGN AOI22FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 14.900 ; # A|0.0@0
      RECT 3.400 13.900 14.800 14.900 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 12.500 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 22.600 7.700 ; # Q|0.0@0
      RECT 21.600 6.700 22.600 17.300 ; # Q|0.0@1
      RECT 6.000 16.300 12.200 17.300 ; # Q|0.0@2
      RECT 19.000 16.300 22.600 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 16.400 11.500 20.000 14.900 ;
      RECT 13.800 16.300 17.400 22.100 ;
      RECT 3.400 18.700 20.000 22.100 ;
    LAYER cont2 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 22.600 5.300 ;
      RECT 6.000 4.300 7.000 7.700 ;
      RECT 16.400 4.300 17.400 7.700 ;
      RECT 0.800 11.500 4.400 12.500 ;
      RECT 8.600 11.500 9.600 12.500 ;
      RECT 13.800 11.500 20.000 12.500 ;
      RECT 6.000 13.900 7.000 22.100 ;
      RECT 16.400 11.500 20.000 14.900 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 13.800 16.300 17.400 22.100 ;
      RECT 0.800 18.700 22.600 19.700 ;
      RECT 0.800 18.700 20.000 22.100 ;
      RECT 0.800 18.700 1.800 24.500 ;
      RECT 11.200 18.700 12.200 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END AOI22FF

MACRO DCFF
  CLASS CORE ;
  FOREIGN DCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 41.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # D|0.0@0
    END
  END D
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 17.300 ; # CN|0.0@0
      RECT 16.400 18.700 17.400 19.700 ; # CN|0.0@1
    END
  END CN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 6.700 40.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.200 9.100 38.200 22.100 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 41.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 41.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 27.800 7.700 ;
      RECT 32.000 6.700 35.600 22.100 ;
      RECT 0.800 9.100 9.600 10.100 ;
      RECT 13.800 6.700 27.800 17.300 ;
      RECT 3.400 9.100 7.000 19.700 ;
      RECT 11.200 11.500 27.800 12.500 ;
      RECT 13.800 13.900 35.600 17.300 ;
      RECT 0.800 16.300 7.000 19.700 ;
      RECT 11.200 16.300 35.600 17.300 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 19.000 13.900 35.600 19.700 ;
      RECT 6.000 18.700 9.600 22.100 ;
      RECT 29.400 13.900 35.600 22.100 ;
      RECT 39.800 21.100 40.800 22.100 ;
    LAYER cont2 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 22.600 0.500 ;
      RECT 29.400 -0.500 33.000 0.500 ;
      RECT 0.800 4.300 25.200 5.300 ;
      RECT 32.000 4.300 35.600 7.700 ;
      RECT 6.000 6.700 27.800 7.700 ;
      RECT 32.000 6.700 40.800 7.700 ;
      RECT 0.800 9.100 4.400 12.500 ;
      RECT 8.600 6.700 27.800 10.100 ;
      RECT 34.600 4.300 35.600 24.500 ;
      RECT 39.800 6.700 40.800 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 4.300 12.200 12.500 ;
      RECT 16.400 6.700 27.800 19.700 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 16.400 13.900 35.600 19.700 ;
      RECT 0.800 16.300 4.400 19.700 ;
      RECT 11.200 16.300 35.600 19.700 ;
      RECT 39.800 16.300 40.800 22.100 ;
      RECT 0.800 18.700 35.600 19.700 ;
      RECT 6.000 18.700 9.600 22.100 ;
      RECT 16.400 4.300 17.400 22.100 ;
      RECT 29.400 13.900 35.600 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 32.000 23.500 38.200 24.500 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
  END
END DCFF

MACRO DCGG
  CLASS CORE ;
  FOREIGN DCGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 49.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # D|0.0@0
    END
  END D
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 17.300 ; # CN|0.0@0
      RECT 11.200 18.700 12.200 19.700 ; # CN|0.0@1
      RECT 32.000 18.700 33.000 22.100 ; # CN|0.0@2
    END
  END CN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 6.700 48.600 17.300 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 6.700 43.400 17.300 ; # QN|0.0@0
      RECT 39.800 18.700 40.800 19.700 ; # QN|0.0@1
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 49.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 49.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 33.000 7.700 ;
      RECT 37.200 6.700 40.800 17.300 ;
      RECT 3.400 9.100 7.000 19.700 ;
      RECT 13.800 9.100 40.800 17.300 ;
      RECT 0.800 16.300 7.000 19.700 ;
      RECT 45.000 16.300 46.000 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 13.800 6.700 17.400 22.100 ;
      RECT 21.600 6.700 30.400 22.100 ;
      RECT 34.600 9.100 38.200 19.700 ;
      RECT 42.400 18.700 48.600 19.700 ;
      RECT 6.000 21.100 30.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 45.000 -0.500 46.000 0.500 ;
      RECT 6.000 4.300 33.000 7.700 ;
      RECT 37.200 4.300 48.600 5.300 ;
      RECT 3.400 6.700 33.000 7.700 ;
      RECT 37.200 4.300 40.800 19.700 ;
      RECT 47.600 4.300 48.600 10.100 ;
      RECT 0.800 9.100 4.400 12.500 ;
      RECT 8.600 4.300 9.600 10.100 ;
      RECT 13.800 9.100 40.800 17.300 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 11.500 40.800 12.500 ;
      RECT 3.400 11.500 7.000 17.300 ;
      RECT 45.000 13.900 46.000 19.700 ;
      RECT 0.800 16.300 7.000 17.300 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 6.000 18.700 9.600 19.700 ;
      RECT 13.800 4.300 17.400 24.500 ;
      RECT 21.600 4.300 30.400 24.500 ;
      RECT 34.600 18.700 48.600 19.700 ;
      RECT 0.800 21.100 4.400 22.100 ;
      RECT 8.600 21.100 30.400 22.100 ;
      RECT 34.600 9.100 35.600 22.100 ;
      RECT 6.000 23.500 9.600 24.500 ;
      RECT 13.800 23.500 33.000 24.500 ;
      RECT 37.200 23.500 38.200 24.500 ;
      RECT 42.400 23.500 43.400 24.500 ;
      RECT 47.600 23.500 48.600 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 20.000 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
  END
END DCGG

MACRO DEC2NDD
  CLASS CORE ;
  FOREIGN DEC2NDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 54.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 9.600 12.500 ; # B|0.0@0
    END
  END B
  PIN EI
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 11.500 20.000 12.500 ; # EI|0.0@0
    END
  END EI
  PIN Q0N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 17.300 ; # Q0N|0.0@0
      RECT 0.800 16.300 7.000 17.300 ; # Q0N|0.0@1
    END
  END Q0N
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 11.500 17.400 12.500 ; # Q1N|0.0@0
      RECT 16.400 16.300 17.400 17.300 ; # Q1N|0.0@1
    END
  END Q1N
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 9.100 53.800 17.300 ; # Q2N|0.0@0
      RECT 50.200 16.300 53.800 17.300 ; # Q2N|0.0@1
    END
  END Q2N
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.200 9.100 38.200 14.900 ; # Q3N|0.0@0
    END
  END Q3N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 54.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 54.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 11.200 6.700 35.600 7.700 ;
      RECT 11.200 6.700 17.400 10.100 ;
      RECT 24.200 6.700 30.400 22.100 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 39.800 9.100 43.400 22.100 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 11.200 6.700 14.800 17.300 ;
      RECT 24.200 11.500 35.600 22.100 ;
      RECT 39.800 11.500 48.600 19.700 ;
      RECT 3.400 13.900 35.600 14.900 ;
      RECT 39.800 13.900 51.200 14.900 ;
      RECT 8.600 13.900 14.800 17.300 ;
      RECT 19.000 13.900 20.000 22.100 ;
      RECT 24.200 16.300 48.600 19.700 ;
      RECT 8.600 13.900 9.600 22.100 ;
      RECT 13.800 18.700 20.000 22.100 ;
      RECT 52.800 18.700 53.800 19.700 ;
      RECT 8.600 21.100 46.000 22.100 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 22.600 0.500 ;
      RECT 32.000 -0.500 35.600 0.500 ;
      RECT 45.000 -0.500 48.600 0.500 ;
      RECT 8.600 4.300 9.600 5.300 ;
      RECT 21.600 4.300 22.600 5.300 ;
      RECT 32.000 4.300 33.000 5.300 ;
      RECT 45.000 4.300 46.000 5.300 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 11.200 6.700 12.200 17.300 ;
      RECT 24.200 6.700 27.800 19.700 ;
      RECT 34.600 6.700 35.600 24.500 ;
      RECT 0.800 9.100 48.600 10.100 ;
      RECT 52.800 9.100 53.800 10.100 ;
      RECT 3.400 9.100 4.400 14.900 ;
      RECT 8.600 9.100 14.800 14.900 ;
      RECT 24.200 9.100 35.600 19.700 ;
      RECT 39.800 9.100 40.800 24.500 ;
      RECT 45.000 11.500 51.200 17.300 ;
      RECT 3.400 13.900 35.600 14.900 ;
      RECT 39.800 13.900 51.200 17.300 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 13.900 7.000 19.700 ;
      RECT 11.200 9.100 14.800 17.300 ;
      RECT 19.000 16.300 53.800 17.300 ;
      RECT 0.800 18.700 7.000 19.700 ;
      RECT 13.800 18.700 48.600 19.700 ;
      RECT 52.800 16.300 53.800 19.700 ;
      RECT 11.200 21.100 22.600 24.500 ;
      RECT 26.800 16.300 46.000 24.500 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 23.500 46.000 24.500 ;
      RECT 50.200 23.500 51.200 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 45.000 28.300 46.000 29.300 ;
      RECT 50.200 28.300 51.200 29.300 ;
  END
END DEC2NDD

MACRO DFFEE
  CLASS CORE ;
  FOREIGN DFFEE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 6.700 30.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 13.900 27.800 22.100 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 24.200 6.700 27.800 12.500 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 16.400 9.100 27.800 12.500 ;
      RECT 3.400 11.500 27.800 12.500 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 11.200 11.500 25.200 17.300 ;
      RECT 6.000 18.700 12.200 22.100 ;
      RECT 16.400 9.100 25.200 22.100 ;
      RECT 3.400 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 30.400 5.300 ;
      RECT 0.800 4.300 20.000 7.700 ;
      RECT 24.200 4.300 30.400 7.700 ;
      RECT 0.800 4.300 1.800 12.500 ;
      RECT 6.000 4.300 12.200 12.500 ;
      RECT 16.400 9.100 27.800 12.500 ;
      RECT 6.000 11.500 27.800 12.500 ;
      RECT 3.400 13.900 7.000 14.900 ;
      RECT 11.200 11.500 25.200 14.900 ;
      RECT 0.800 16.300 4.400 17.300 ;
      RECT 13.800 11.500 25.200 22.100 ;
      RECT 29.400 16.300 30.400 22.100 ;
      RECT 8.600 18.700 25.200 22.100 ;
      RECT 0.800 21.100 4.400 24.500 ;
      RECT 0.800 23.500 7.000 24.500 ;
      RECT 11.200 18.700 14.800 24.500 ;
      RECT 21.600 23.500 27.800 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END DFFEE

MACRO DFFFF
  CLASS CORE ;
  FOREIGN DFFFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 33.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 6.700 33.000 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 6.700 30.400 22.100 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 33.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 33.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 27.800 7.700 ;
      RECT 0.800 9.100 14.800 10.100 ;
      RECT 19.000 6.700 27.800 19.700 ;
      RECT 3.400 11.500 27.800 12.500 ;
      RECT 3.400 9.100 7.000 22.100 ;
      RECT 11.200 11.500 27.800 19.700 ;
      RECT 3.400 21.100 14.800 22.100 ;
      RECT 19.000 6.700 22.600 22.100 ;
      RECT 26.800 6.700 27.800 22.100 ;
      RECT 32.000 21.100 33.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 33.000 5.300 ;
      RECT 6.000 6.700 27.800 10.100 ;
      RECT 32.000 4.300 33.000 10.100 ;
      RECT 0.800 9.100 27.800 10.100 ;
      RECT 0.800 9.100 17.400 12.500 ;
      RECT 21.600 4.300 27.800 14.900 ;
      RECT 3.400 9.100 7.000 14.900 ;
      RECT 11.200 13.900 27.800 14.900 ;
      RECT 3.400 9.100 4.400 24.500 ;
      RECT 11.200 13.900 20.000 19.700 ;
      RECT 24.200 4.300 27.800 22.100 ;
      RECT 32.000 16.300 33.000 22.100 ;
      RECT 3.400 18.700 7.000 24.500 ;
      RECT 3.400 21.100 14.800 24.500 ;
      RECT 19.000 21.100 27.800 22.100 ;
      RECT 0.800 23.500 14.800 24.500 ;
      RECT 19.000 21.100 22.600 24.500 ;
      RECT 26.800 23.500 30.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 12.200 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
  END
END DFFFF

MACRO DFFGG
  CLASS CORE ;
  FOREIGN DFFGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 41.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 6.700 40.800 14.900 ; # Q|0.0@0
      RECT 37.200 13.900 40.800 14.900 ; # Q|0.0@1
      RECT 37.200 13.900 38.200 19.700 ; # Q|0.0@2
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 6.700 35.600 17.300 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 41.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 41.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 6.000 6.700 27.800 10.100 ;
      RECT 32.000 6.700 33.000 22.100 ;
      RECT 0.800 9.100 27.800 10.100 ;
      RECT 3.400 9.100 7.000 22.100 ;
      RECT 11.200 11.500 33.000 14.900 ;
      RECT 3.400 13.900 33.000 14.900 ;
      RECT 3.400 13.900 14.800 22.100 ;
      RECT 19.000 11.500 33.000 19.700 ;
      RECT 3.400 18.700 33.000 19.700 ;
      RECT 3.400 18.700 27.800 22.100 ;
      RECT 37.200 21.100 38.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 6.000 4.300 22.600 5.300 ;
      RECT 26.800 4.300 35.600 7.700 ;
      RECT 39.800 4.300 40.800 10.100 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 24.200 6.700 35.600 7.700 ;
      RECT 0.800 6.700 1.800 12.500 ;
      RECT 8.600 9.100 30.400 10.100 ;
      RECT 34.600 4.300 35.600 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 9.100 25.200 12.500 ;
      RECT 29.400 4.300 30.400 24.500 ;
      RECT 37.200 11.500 38.200 12.500 ;
      RECT 3.400 13.900 17.400 14.900 ;
      RECT 21.600 13.900 33.000 14.900 ;
      RECT 0.800 16.300 12.200 17.300 ;
      RECT 19.000 16.300 22.600 24.500 ;
      RECT 26.800 13.900 33.000 22.100 ;
      RECT 37.200 16.300 40.800 22.100 ;
      RECT 0.800 16.300 7.000 22.100 ;
      RECT 11.200 18.700 22.600 19.700 ;
      RECT 26.800 18.700 40.800 22.100 ;
      RECT 16.400 18.700 22.600 24.500 ;
      RECT 3.400 23.500 30.400 24.500 ;
      RECT 34.600 18.700 35.600 24.500 ;
      RECT 39.800 16.300 40.800 24.500 ;
      RECT 0.800 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
  END
END DFFGG

MACRO DPCFF
  CLASS CORE ;
  FOREIGN DPCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 54.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 13.900 40.800 17.300 ; # PN|0.0@0
      RECT 37.200 16.300 40.800 17.300 ; # PN|0.0@1
    END
  END PN
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 13.900 38.200 14.900 ; # CN|0.0@0
    END
  END CN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 6.700 53.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 11.500 48.600 22.100 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 54.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 54.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 51.200 10.100 ;
      RECT 0.800 9.100 51.200 10.100 ;
      RECT 3.400 6.700 46.000 12.500 ;
      RECT 50.200 6.700 51.200 14.900 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 13.800 6.700 33.000 14.900 ;
      RECT 42.400 6.700 46.000 22.100 ;
      RECT 13.800 6.700 14.800 22.100 ;
      RECT 19.000 6.700 33.000 22.100 ;
      RECT 3.400 18.700 33.000 22.100 ;
      RECT 37.200 18.700 46.000 22.100 ;
      RECT 3.400 21.100 46.000 22.100 ;
      RECT 52.800 21.100 53.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 16.400 -0.500 22.600 0.500 ;
      RECT 50.200 -0.500 51.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 27.800 7.700 ;
      RECT 32.000 4.300 51.200 5.300 ;
      RECT 6.000 6.700 27.800 7.700 ;
      RECT 32.000 4.300 35.600 17.300 ;
      RECT 39.800 4.300 48.600 10.100 ;
      RECT 52.800 6.700 53.800 10.100 ;
      RECT 0.800 9.100 9.600 12.500 ;
      RECT 13.800 9.100 48.600 10.100 ;
      RECT 0.800 11.500 46.000 12.500 ;
      RECT 50.200 11.500 51.200 14.900 ;
      RECT 3.400 9.100 7.000 24.500 ;
      RECT 11.200 11.500 35.600 14.900 ;
      RECT 42.400 4.300 46.000 14.900 ;
      RECT 13.800 16.300 38.200 17.300 ;
      RECT 45.000 4.300 46.000 24.500 ;
      RECT 52.800 16.300 53.800 22.100 ;
      RECT 3.400 18.700 33.000 24.500 ;
      RECT 37.200 18.700 48.600 24.500 ;
      RECT 3.400 21.100 48.600 24.500 ;
      RECT 0.800 23.500 51.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
      RECT 50.200 28.300 51.200 29.300 ;
  END
END DPCFF

MACRO DPFF
  CLASS CORE ;
  FOREIGN DPFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 44.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 9.100 33.000 14.900 ; # PN|0.0@0
    END
  END PN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 6.700 43.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.200 9.100 38.200 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 44.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 44.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 38.200 7.700 ;
      RECT 3.400 9.100 14.800 12.500 ;
      RECT 19.000 6.700 30.400 19.700 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 3.400 11.500 30.400 12.500 ;
      RECT 3.400 9.100 7.000 22.100 ;
      RECT 13.800 11.500 30.400 19.700 ;
      RECT 13.800 16.300 35.600 19.700 ;
      RECT 3.400 21.100 27.800 22.100 ;
      RECT 34.600 21.100 38.200 22.100 ;
      RECT 42.400 21.100 43.400 22.100 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 37.200 -0.500 40.800 0.500 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 16.400 4.300 17.400 5.300 ;
      RECT 21.600 4.300 25.200 7.700 ;
      RECT 29.400 4.300 38.200 7.700 ;
      RECT 3.400 6.700 9.600 12.500 ;
      RECT 19.000 6.700 38.200 7.700 ;
      RECT 42.400 6.700 43.400 10.100 ;
      RECT 0.800 9.100 14.800 12.500 ;
      RECT 19.000 6.700 22.600 14.900 ;
      RECT 26.800 6.700 27.800 22.100 ;
      RECT 34.600 4.300 38.200 10.100 ;
      RECT 0.800 11.500 30.400 12.500 ;
      RECT 3.400 6.700 7.000 14.900 ;
      RECT 13.800 11.500 30.400 14.900 ;
      RECT 0.800 16.300 4.400 24.500 ;
      RECT 13.800 11.500 17.400 24.500 ;
      RECT 21.600 16.300 33.000 19.700 ;
      RECT 42.400 16.300 43.400 22.100 ;
      RECT 0.800 18.700 7.000 24.500 ;
      RECT 13.800 18.700 35.600 19.700 ;
      RECT 0.800 21.100 17.400 24.500 ;
      RECT 21.600 11.500 30.400 22.100 ;
      RECT 34.600 21.100 38.200 22.100 ;
      RECT 0.800 23.500 25.200 24.500 ;
      RECT 29.400 11.500 30.400 24.500 ;
      RECT 34.600 18.700 35.600 24.500 ;
      RECT 39.800 23.500 40.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 26.800 28.300 30.400 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
  END
END DPFF

MACRO INVDD
  CLASS CORE ;
  FOREIGN INVDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 3.400 9.100 4.400 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 28.300 4.400 29.300 ;
  END
END INVDD

MACRO INVFF
  CLASS CORE ;
  FOREIGN INVFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 19.700 ; # Q|0.0@0
      RECT 0.800 18.700 4.400 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 21.100 4.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 0.800 9.100 4.400 10.100 ;
      RECT 3.400 9.100 4.400 12.500 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 0.800 21.100 4.400 22.100 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END INVFF

MACRO INVGG
  CLASS CORE ;
  FOREIGN INVGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 6.000 6.700 7.000 12.500 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END INVGG

MACRO INVHH
  CLASS CORE ;
  FOREIGN INVHH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 7.000 5.300 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END INVHH

MACRO INVII
  CLASS CORE ;
  FOREIGN INVII 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # Q|0.0@0
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@1
      RECT 3.400 16.300 9.600 17.300 ; # Q|0.0@2
      RECT 3.400 16.300 4.400 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 5.700 21.600 7.300 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 3.400 11.500 7.000 12.500 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 6.000 21.100 7.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 9.600 5.300 ;
      RECT 3.400 4.300 7.000 14.900 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 3.400 4.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 6.000 18.700 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END INVII

MACRO INVJJ
  CLASS CORE ;
  FOREIGN INVJJ 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 19.700 ; # Q|0.0@0
      RECT 8.600 6.700 9.600 14.900 ; # Q|0.0@1
      RECT 13.800 16.300 14.800 19.700 ; # Q|0.0@2
      RECT 3.400 18.700 14.800 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ;
      RECT 13.800 13.900 14.800 14.900 ;
      RECT 6.000 16.300 12.200 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 7.000 5.300 ;
      RECT 11.200 4.300 12.200 5.300 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 8.600 6.700 9.600 10.100 ;
      RECT 3.400 9.100 9.600 10.100 ;
      RECT 6.000 9.100 7.000 12.500 ;
      RECT 13.800 13.900 14.800 19.700 ;
      RECT 3.400 16.300 14.800 17.300 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END INVJJ

MACRO INVJK
  CLASS CORE ;
  FOREIGN INVJK 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 17.400 12.500 ; # A|0.0@0
      RECT 16.400 11.500 17.400 14.900 ; # A|0.0@1
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 12.200 10.100 ; # Q|0.0@0
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@1
      RECT 8.600 9.100 9.600 14.900 ; # Q|0.0@2
      RECT 13.800 16.300 14.800 19.700 ; # Q|0.0@3
      RECT 3.400 18.700 14.800 19.700 ; # Q|0.0@4
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 11.200 6.700 14.800 7.700 ;
      RECT 13.800 6.700 14.800 10.100 ;
      RECT 13.800 13.900 14.800 14.900 ;
      RECT 6.000 16.300 12.200 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 16.400 4.300 17.400 5.300 ;
      RECT 3.400 6.700 14.800 7.700 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 11.200 6.700 14.800 12.500 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 11.200 11.500 17.400 12.500 ;
      RECT 13.800 6.700 14.800 19.700 ;
      RECT 3.400 16.300 14.800 17.300 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END INVJK

MACRO INVKK
  CLASS CORE ;
  FOREIGN INVKK 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 20.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 6.700 20.000 19.700 ; # Q|0.0@0
      RECT 8.600 9.100 20.000 10.100 ; # Q|0.0@1
      RECT 3.400 16.300 4.400 19.700 ; # Q|0.0@2
      RECT 3.400 18.700 20.000 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 20.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 20.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 14.900 ;
      RECT 11.200 6.700 14.800 7.700 ;
      RECT 3.400 13.900 9.600 14.900 ;
      RECT 13.800 13.900 14.800 17.300 ;
      RECT 6.000 16.300 17.400 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 13.800 4.300 17.400 7.700 ;
      RECT 3.400 6.700 20.000 7.700 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 11.200 6.700 12.200 12.500 ;
      RECT 19.000 6.700 20.000 10.100 ;
      RECT 0.800 11.500 17.400 12.500 ;
      RECT 3.400 11.500 9.600 17.300 ;
      RECT 13.800 11.500 14.800 19.700 ;
      RECT 3.400 16.300 20.000 17.300 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 11.500 9.600 19.700 ;
      RECT 19.000 16.300 20.000 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END INVKK

MACRO JKCFF
  CLASS CORE ;
  FOREIGN JKCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 52.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 11.500 40.800 12.500 ; # CN|0.0@0
    END
  END CN
  PIN JN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # JN|0.0@0
    END
  END JN
  PIN K
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # K|0.0@0
    END
  END K
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 50.200 6.700 51.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 9.100 48.600 22.100 ; # QN|0.0@0
      RECT 0.800 16.300 1.800 22.100 ; # QN|0.0@1
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 52.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 52.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 33.000 10.100 ;
      RECT 42.400 6.700 48.600 7.700 ;
      RECT 6.000 9.100 46.000 10.100 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 8.600 9.100 38.200 12.500 ;
      RECT 42.400 6.700 46.000 22.100 ;
      RECT 8.600 6.700 9.600 22.100 ;
      RECT 13.800 13.900 46.000 17.300 ;
      RECT 6.000 16.300 9.600 22.100 ;
      RECT 3.400 18.700 22.600 22.100 ;
      RECT 32.000 13.900 46.000 22.100 ;
      RECT 3.400 21.100 46.000 22.100 ;
      RECT 50.200 21.100 51.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 9.600 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 26.800 -0.500 27.800 0.500 ;
      RECT 39.800 -0.500 43.400 0.500 ;
      RECT 47.600 -0.500 48.600 0.500 ;
      RECT 0.800 4.300 33.000 5.300 ;
      RECT 42.400 4.300 51.200 7.700 ;
      RECT 6.000 6.700 51.200 7.700 ;
      RECT 6.000 6.700 38.200 10.100 ;
      RECT 42.400 4.300 46.000 24.500 ;
      RECT 50.200 4.300 51.200 10.100 ;
      RECT 0.800 11.500 4.400 12.500 ;
      RECT 11.200 6.700 38.200 12.500 ;
      RECT 0.800 11.500 1.800 19.700 ;
      RECT 13.800 13.900 46.000 24.500 ;
      RECT 0.800 16.300 7.000 19.700 ;
      RECT 11.200 16.300 46.000 24.500 ;
      RECT 50.200 16.300 51.200 22.100 ;
      RECT 0.800 18.700 46.000 19.700 ;
      RECT 3.400 18.700 46.000 24.500 ;
      RECT 0.800 23.500 48.600 24.500 ;
      RECT 0.800 28.300 9.600 29.300 ;
      RECT 13.800 28.300 17.400 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
  END
END JKCFF

MACRO JKCGG
  CLASS CORE ;
  FOREIGN JKCGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 59.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 10.100 ; # CN|0.0@0
      RECT 32.000 18.700 33.000 19.700 ; # CN|0.0@1
    END
  END CN
  PIN JN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 13.900 56.400 14.900 ; # JN|0.0@0
    END
  END JN
  PIN K
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 50.200 11.500 51.200 14.900 ; # K|0.0@0
    END
  END K
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 6.700 56.400 7.700 ; # Q|0.0@0
      RECT 47.600 9.100 48.600 10.100 ; # Q|0.0@1
      RECT 58.000 9.100 59.000 12.500 ; # Q|0.0@2
      RECT 45.000 11.500 46.000 14.900 ; # Q|0.0@3
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 6.700 43.400 7.700 ; # QN|0.0@0
      RECT 42.400 11.500 43.400 19.700 ; # QN|0.0@1
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 59.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 59.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 6.000 6.700 27.800 7.700 ;
      RECT 37.200 6.700 38.200 22.100 ;
      RECT 45.000 6.700 53.800 7.700 ;
      RECT 58.000 6.700 59.000 7.700 ;
      RECT 0.800 9.100 7.000 10.100 ;
      RECT 13.800 9.100 46.000 10.100 ;
      RECT 50.200 6.700 53.800 10.100 ;
      RECT 3.400 11.500 22.600 14.900 ;
      RECT 26.800 9.100 40.800 14.900 ;
      RECT 52.800 11.500 56.400 12.500 ;
      RECT 3.400 13.900 40.800 14.900 ;
      RECT 52.800 6.700 53.800 22.100 ;
      RECT 58.000 13.900 59.000 14.900 ;
      RECT 3.400 11.500 17.400 19.700 ;
      RECT 21.600 13.900 27.800 22.100 ;
      RECT 32.000 9.100 40.800 17.300 ;
      RECT 45.000 16.300 56.400 22.100 ;
      RECT 0.800 18.700 30.400 19.700 ;
      RECT 34.600 9.100 40.800 22.100 ;
      RECT 0.800 18.700 1.800 22.100 ;
      RECT 6.000 21.100 56.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 50.200 -0.500 51.200 0.500 ;
      RECT 58.000 -0.500 59.000 0.500 ;
      RECT 6.000 4.300 27.800 7.700 ;
      RECT 32.000 4.300 33.000 5.300 ;
      RECT 37.200 4.300 46.000 5.300 ;
      RECT 0.800 6.700 1.800 12.500 ;
      RECT 34.600 6.700 38.200 24.500 ;
      RECT 42.400 6.700 53.800 10.100 ;
      RECT 58.000 6.700 59.000 7.700 ;
      RECT 11.200 9.100 56.400 10.100 ;
      RECT 0.800 11.500 40.800 12.500 ;
      RECT 52.800 11.500 59.000 12.500 ;
      RECT 3.400 11.500 40.800 14.900 ;
      RECT 47.600 13.900 51.200 24.500 ;
      RECT 58.000 11.500 59.000 14.900 ;
      RECT 8.600 11.500 17.400 24.500 ;
      RECT 21.600 9.100 40.800 17.300 ;
      RECT 45.000 16.300 56.400 24.500 ;
      RECT 0.800 18.700 1.800 22.100 ;
      RECT 6.000 18.700 30.400 24.500 ;
      RECT 34.600 9.100 40.800 24.500 ;
      RECT 6.000 21.100 56.400 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 29.400 28.300 33.000 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 55.400 28.300 59.000 29.300 ;
  END
END JKCGG

MACRO JKPCFF
  CLASS CORE ;
  FOREIGN JKPCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 70.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 11.500 43.400 14.900 ; # PN|0.0@0
    END
  END PN
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.200 16.300 38.200 17.300 ; # CN|0.0@0
    END
  END CN
  PIN JN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 63.200 13.900 64.200 14.900 ; # JN|0.0@0
    END
  END JN
  PIN K
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 68.400 11.500 69.400 14.900 ; # K|0.0@0
    END
  END K
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 58.000 13.900 59.000 14.900 ; # Q|0.0@0
      RECT 58.000 18.700 59.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 9.100 56.400 17.300 ; # QN|0.0@0
      RECT 60.600 18.700 61.600 22.100 ; # QN|0.0@1
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 70.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 70.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 66.800 7.700 ;
      RECT 3.400 6.700 25.200 22.100 ;
      RECT 29.400 6.700 53.800 10.100 ;
      RECT 58.000 6.700 66.800 10.100 ;
      RECT 29.400 6.700 40.800 14.900 ;
      RECT 45.000 6.700 53.800 22.100 ;
      RECT 58.000 6.700 61.600 12.500 ;
      RECT 65.800 6.700 66.800 22.100 ;
      RECT 60.600 6.700 61.600 17.300 ;
      RECT 3.400 16.300 35.600 22.100 ;
      RECT 39.800 16.300 53.800 17.300 ;
      RECT 58.000 16.300 69.400 17.300 ;
      RECT 3.400 18.700 38.200 22.100 ;
      RECT 42.400 18.700 56.400 22.100 ;
      RECT 63.200 16.300 69.400 22.100 ;
      RECT 3.400 21.100 59.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 52.800 -0.500 53.800 0.500 ;
      RECT 58.000 -0.500 66.800 0.500 ;
      RECT 0.800 4.300 66.800 5.300 ;
      RECT 6.000 4.300 66.800 7.700 ;
      RECT 0.800 9.100 25.200 12.500 ;
      RECT 29.400 4.300 30.400 12.500 ;
      RECT 34.600 4.300 53.800 10.100 ;
      RECT 58.000 4.300 66.800 10.100 ;
      RECT 29.400 11.500 40.800 12.500 ;
      RECT 45.000 4.300 53.800 17.300 ;
      RECT 58.000 4.300 61.600 12.500 ;
      RECT 3.400 9.100 4.400 24.500 ;
      RECT 8.600 4.300 25.200 14.900 ;
      RECT 32.000 11.500 40.800 14.900 ;
      RECT 60.600 4.300 61.600 17.300 ;
      RECT 68.400 13.900 69.400 24.500 ;
      RECT 8.600 4.300 22.600 24.500 ;
      RECT 26.800 16.300 35.600 17.300 ;
      RECT 39.800 16.300 53.800 17.300 ;
      RECT 58.000 16.300 69.400 17.300 ;
      RECT 3.400 18.700 25.200 24.500 ;
      RECT 29.400 18.700 43.400 24.500 ;
      RECT 47.600 18.700 56.400 24.500 ;
      RECT 63.200 16.300 69.400 24.500 ;
      RECT 3.400 21.100 59.000 24.500 ;
      RECT 0.800 23.500 69.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 52.800 28.300 56.400 29.300 ;
      RECT 60.600 28.300 69.400 29.300 ;
  END
END JKPCFF

MACRO JKPCGG
  CLASS CORE ;
  FOREIGN JKPCGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 88.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 63.200 11.500 64.200 12.500 ; # PN|0.0@0
    END
  END PN
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 71.000 6.700 72.000 10.100 ; # CN|0.0@0
      RECT 24.200 9.100 25.200 12.500 ; # CN|0.0@1
    END
  END CN
  PIN JN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # JN|0.0@0
    END
  END JN
  PIN K
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # K|0.0@0
    END
  END K
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 78.800 11.500 79.800 22.100 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 86.600 6.700 87.600 7.700 ; # QN|0.0@0
      RECT 8.600 11.500 9.600 22.100 ; # QN|0.0@1
      RECT 84.000 11.500 85.000 22.100 ; # QN|0.0@2
      RECT 0.800 16.300 1.800 22.100 ; # QN|0.0@3
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 88.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 88.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 69.400 7.700 ;
      RECT 73.600 6.700 85.000 10.100 ;
      RECT 3.400 6.700 22.600 10.100 ;
      RECT 26.800 6.700 48.600 14.900 ;
      RECT 52.800 6.700 64.200 10.100 ;
      RECT 73.600 9.100 87.600 10.100 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 13.800 6.700 22.600 17.300 ;
      RECT 26.800 11.500 61.600 14.900 ;
      RECT 65.800 11.500 77.200 22.100 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 13.800 13.900 77.200 14.900 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 11.200 16.300 40.800 17.300 ;
      RECT 45.000 13.900 77.200 22.100 ;
      RECT 11.200 16.300 20.000 22.100 ;
      RECT 26.800 18.700 77.200 22.100 ;
      RECT 11.200 21.100 77.200 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 14.800 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 39.800 -0.500 40.800 0.500 ;
      RECT 68.400 -0.500 72.000 0.500 ;
      RECT 76.200 -0.500 77.200 0.500 ;
      RECT 81.400 -0.500 82.400 0.500 ;
      RECT 3.400 4.300 87.600 5.300 ;
      RECT 3.400 4.300 69.400 7.700 ;
      RECT 73.600 4.300 87.600 10.100 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 6.000 4.300 22.600 10.100 ;
      RECT 26.800 4.300 48.600 14.900 ;
      RECT 52.800 4.300 64.200 10.100 ;
      RECT 71.000 9.100 87.600 10.100 ;
      RECT 13.800 4.300 22.600 17.300 ;
      RECT 26.800 11.500 61.600 14.900 ;
      RECT 65.800 11.500 77.200 24.500 ;
      RECT 0.800 13.900 1.800 17.300 ;
      RECT 13.800 13.900 77.200 14.900 ;
      RECT 6.000 16.300 7.000 24.500 ;
      RECT 11.200 16.300 40.800 17.300 ;
      RECT 45.000 13.900 77.200 24.500 ;
      RECT 3.400 18.700 7.000 24.500 ;
      RECT 11.200 16.300 20.000 22.100 ;
      RECT 26.800 18.700 79.800 24.500 ;
      RECT 84.000 18.700 85.000 24.500 ;
      RECT 11.200 21.100 79.800 22.100 ;
      RECT 0.800 23.500 9.600 24.500 ;
      RECT 13.800 4.300 14.800 24.500 ;
      RECT 19.000 21.100 79.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
      RECT 50.200 28.300 51.200 29.300 ;
      RECT 63.200 28.300 64.200 29.300 ;
      RECT 68.400 28.300 69.400 29.300 ;
      RECT 76.200 28.300 77.200 29.300 ;
      RECT 81.400 28.300 82.400 29.300 ;
      RECT 86.600 28.300 87.600 29.300 ;
  END
END JKPCGG

MACRO JKPCHH
  CLASS CORE ;
  FOREIGN JKPCHH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 93.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 16.300 12.200 17.300 ; # CLK|0.0@0
    END
  END CLK
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 58.000 9.100 59.000 10.100 ; # PN|0.0@0
    END
  END PN
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 25.200 12.500 ; # CN|0.0@0
      RECT 68.400 18.700 69.400 19.700 ; # CN|0.0@1
    END
  END CN
  PIN JN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # JN|0.0@0
    END
  END JN
  PIN K
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # K|0.0@0
    END
  END K
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 84.000 6.700 85.000 10.100 ; # Q|0.0@0
      RECT 86.600 11.500 87.600 22.100 ; # Q|0.0@1
      RECT 84.000 18.700 87.600 22.100 ; # Q|0.0@2
      RECT 76.200 21.100 87.600 22.100 ; # Q|0.0@3
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 89.200 6.700 92.800 7.700 ; # QN|0.0@0
      RECT 89.200 6.700 90.200 14.900 ; # QN|0.0@1
      RECT 8.600 11.500 12.200 12.500 ; # QN|0.0@2
      RECT 8.600 16.300 9.600 22.100 ; # QN|0.0@3
      RECT 89.200 18.700 90.200 19.700 ; # QN|0.0@4
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 93.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 93.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 69.400 7.700 ;
      RECT 73.600 6.700 77.200 10.100 ;
      RECT 81.400 6.700 82.400 17.300 ;
      RECT 86.600 6.700 87.600 10.100 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 13.800 6.700 56.400 10.100 ;
      RECT 63.200 9.100 82.400 10.100 ;
      RECT 13.800 6.700 20.000 22.100 ;
      RECT 26.800 11.500 59.000 12.500 ;
      RECT 63.200 9.100 72.000 17.300 ;
      RECT 76.200 11.500 85.000 17.300 ;
      RECT 91.800 11.500 92.800 19.700 ;
      RECT 0.800 13.900 4.400 22.100 ;
      RECT 8.600 13.900 30.400 14.900 ;
      RECT 39.800 13.900 85.000 17.300 ;
      RECT 13.800 13.900 30.400 17.300 ;
      RECT 37.200 16.300 85.000 17.300 ;
      RECT 89.200 16.300 92.800 17.300 ;
      RECT 0.800 18.700 7.000 22.100 ;
      RECT 26.800 18.700 66.800 19.700 ;
      RECT 71.000 13.900 79.800 19.700 ;
      RECT 13.800 21.100 43.400 22.100 ;
      RECT 47.600 21.100 74.600 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 17.400 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 55.400 -0.500 59.000 0.500 ;
      RECT 71.000 -0.500 72.000 0.500 ;
      RECT 84.000 -0.500 85.000 0.500 ;
      RECT 89.200 -0.500 90.200 0.500 ;
      RECT 6.000 4.300 72.000 7.700 ;
      RECT 78.800 4.300 92.800 5.300 ;
      RECT 3.400 6.700 82.400 7.700 ;
      RECT 86.600 4.300 87.600 10.100 ;
      RECT 91.800 4.300 92.800 7.700 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 8.600 4.300 48.600 10.100 ;
      RECT 52.800 4.300 59.000 24.500 ;
      RECT 63.200 4.300 69.400 17.300 ;
      RECT 78.800 4.300 82.400 12.500 ;
      RECT 3.400 11.500 4.400 24.500 ;
      RECT 11.200 4.300 20.000 14.900 ;
      RECT 26.800 11.500 59.000 12.500 ;
      RECT 63.200 11.500 74.600 17.300 ;
      RECT 78.800 11.500 85.000 12.500 ;
      RECT 91.800 11.500 92.800 19.700 ;
      RECT 0.800 13.900 30.400 14.900 ;
      RECT 39.800 13.900 79.800 17.300 ;
      RECT 84.000 11.500 85.000 19.700 ;
      RECT 0.800 13.900 4.400 24.500 ;
      RECT 13.800 4.300 17.400 24.500 ;
      RECT 24.200 16.300 85.000 17.300 ;
      RECT 89.200 16.300 92.800 19.700 ;
      RECT 0.800 18.700 7.000 24.500 ;
      RECT 11.200 18.700 20.000 22.100 ;
      RECT 26.800 16.300 66.800 24.500 ;
      RECT 71.000 13.900 79.800 19.700 ;
      RECT 11.200 21.100 74.600 22.100 ;
      RECT 89.200 16.300 90.200 22.100 ;
      RECT 0.800 23.500 17.400 24.500 ;
      RECT 21.600 23.500 77.200 24.500 ;
      RECT 81.400 23.500 82.400 24.500 ;
      RECT 86.600 23.500 87.600 24.500 ;
      RECT 91.800 23.500 92.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 22.600 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 52.800 28.300 56.400 29.300 ;
      RECT 71.000 28.300 72.000 29.300 ;
      RECT 76.200 28.300 77.200 29.300 ;
      RECT 81.400 28.300 82.400 29.300 ;
      RECT 86.600 28.300 87.600 29.300 ;
      RECT 91.800 28.300 92.800 29.300 ;
  END
END JKPCHH

MACRO KEEP
  CLASS CORE ;
  FOREIGN KEEP 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN DBUS
    DIRECTION INOUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # DBUS|0.0@0
    END
  END DBUS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 0.800 21.100 4.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 4.300 7.000 5.300 ;
      RECT 3.400 4.300 7.000 17.300 ;
      RECT 0.800 11.500 7.000 14.900 ;
      RECT 3.400 4.300 4.400 22.100 ;
      RECT 0.800 21.100 4.400 22.100 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
  END
END KEEP

MACRO LTCFF
  CLASS CORE ;
  FOREIGN LTCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 16.300 9.600 17.300 ; # D|0.0@0
    END
  END D
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 19.700 ; # CN|0.0@0
    END
  END CN
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # S|0.0@0
    END
  END S
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 17.300 ; # Q|0.0@0
      RECT 21.600 16.300 25.200 17.300 ; # Q|0.0@1
      RECT 21.600 16.300 22.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 6.700 27.800 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 21.600 6.700 22.600 14.900 ;
      RECT 3.400 9.100 22.600 10.100 ;
      RECT 3.400 6.700 9.600 14.900 ;
      RECT 13.800 9.100 22.600 14.900 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 13.800 9.100 20.000 22.100 ;
      RECT 6.000 6.700 7.000 22.100 ;
      RECT 3.400 21.100 7.000 22.100 ;
      RECT 26.800 21.100 27.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 9.600 0.500 ;
      RECT 21.600 -0.500 25.200 0.500 ;
      RECT 0.800 4.300 25.200 5.300 ;
      RECT 3.400 4.300 22.600 10.100 ;
      RECT 26.800 6.700 27.800 10.100 ;
      RECT 3.400 4.300 9.600 14.900 ;
      RECT 13.800 4.300 22.600 14.900 ;
      RECT 0.800 13.900 9.600 14.900 ;
      RECT 0.800 13.900 4.400 17.300 ;
      RECT 13.800 4.300 17.400 24.500 ;
      RECT 26.800 16.300 27.800 22.100 ;
      RECT 3.400 18.700 7.000 22.100 ;
      RECT 11.200 18.700 17.400 22.100 ;
      RECT 21.600 18.700 27.800 19.700 ;
      RECT 0.800 21.100 7.000 22.100 ;
      RECT 11.200 21.100 22.600 22.100 ;
      RECT 0.800 21.100 4.400 24.500 ;
      RECT 13.800 21.100 20.000 24.500 ;
      RECT 24.200 23.500 25.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 17.400 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END LTCFF

MACRO LTCGG
  CLASS CORE ;
  FOREIGN LTCGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 36.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 16.300 9.600 17.300 ; # D|0.0@0
    END
  END D
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 11.500 20.000 12.500 ; # CN|0.0@0
    END
  END CN
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # S|0.0@0
    END
  END S
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 6.700 30.400 17.300 ; # Q|0.0@0
      RECT 26.800 18.700 27.800 19.700 ; # Q|0.0@1
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 6.700 35.600 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 36.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 36.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 4.400 7.700 ;
      RECT 8.600 6.700 27.800 10.100 ;
      RECT 3.400 9.100 27.800 10.100 ;
      RECT 3.400 9.100 17.400 14.900 ;
      RECT 21.600 6.700 27.800 17.300 ;
      RECT 3.400 13.900 27.800 14.900 ;
      RECT 32.000 13.900 33.000 19.700 ;
      RECT 3.400 9.100 7.000 19.700 ;
      RECT 11.200 13.900 27.800 17.300 ;
      RECT 11.200 6.700 17.400 22.100 ;
      RECT 21.600 6.700 25.200 19.700 ;
      RECT 29.400 18.700 33.000 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 0.800 4.300 7.000 5.300 ;
      RECT 13.800 4.300 17.400 22.100 ;
      RECT 21.600 4.300 35.600 5.300 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 8.600 6.700 27.800 10.100 ;
      RECT 34.600 4.300 35.600 10.100 ;
      RECT 6.000 9.100 27.800 10.100 ;
      RECT 0.800 11.500 17.400 12.500 ;
      RECT 21.600 4.300 27.800 19.700 ;
      RECT 3.400 13.900 27.800 14.900 ;
      RECT 32.000 13.900 33.000 19.700 ;
      RECT 3.400 11.500 7.000 22.100 ;
      RECT 11.200 13.900 27.800 17.300 ;
      RECT 11.200 6.700 17.400 22.100 ;
      RECT 21.600 18.700 33.000 19.700 ;
      RECT 0.800 23.500 4.400 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 29.400 23.500 30.400 24.500 ;
      RECT 34.600 23.500 35.600 24.500 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 19.000 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
  END
END LTCGG

MACRO LTFF
  CLASS CORE ;
  FOREIGN LTFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # S|0.0@0
    END
  END S
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 6.700 22.600 19.700 ; # Q|0.0@0
      RECT 19.000 18.700 22.600 19.700 ; # Q|0.0@1
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 11.200 6.700 20.000 14.900 ;
      RECT 3.400 9.100 20.000 10.100 ;
      RECT 11.200 6.700 12.200 22.100 ;
      RECT 16.400 6.700 20.000 17.300 ;
      RECT 6.000 6.700 7.000 22.100 ;
      RECT 16.400 6.700 17.400 22.100 ;
      RECT 3.400 21.100 7.000 22.100 ;
      RECT 24.200 21.100 25.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 16.400 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 7.000 5.300 ;
      RECT 11.200 4.300 22.600 5.300 ;
      RECT 3.400 4.300 7.000 14.900 ;
      RECT 11.200 4.300 20.000 14.900 ;
      RECT 24.200 6.700 25.200 10.100 ;
      RECT 0.800 9.100 7.000 12.500 ;
      RECT 3.400 13.900 20.000 14.900 ;
      RECT 0.800 16.300 4.400 24.500 ;
      RECT 11.200 4.300 14.800 17.300 ;
      RECT 19.000 4.300 20.000 19.700 ;
      RECT 24.200 16.300 25.200 22.100 ;
      RECT 0.800 18.700 7.000 22.100 ;
      RECT 11.200 4.300 12.200 22.100 ;
      RECT 16.400 18.700 20.000 19.700 ;
      RECT 16.400 18.700 17.400 24.500 ;
      RECT 13.800 23.500 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END LTFF

MACRO LTGG
  CLASS CORE ;
  FOREIGN LTGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # S|0.0@0
    END
  END S
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 17.300 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 6.700 30.400 17.300 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 21.600 6.700 22.600 19.700 ;
      RECT 3.400 9.100 22.600 12.500 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 11.200 9.100 22.600 17.300 ;
      RECT 26.800 13.900 27.800 19.700 ;
      RECT 0.800 18.700 7.000 19.700 ;
      RECT 13.800 6.700 14.800 22.100 ;
      RECT 19.000 18.700 30.400 19.700 ;
      RECT 0.800 18.700 1.800 22.100 ;
      RECT 6.000 6.700 7.000 22.100 ;
      RECT 11.200 21.100 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 16.400 -0.500 22.600 0.500 ;
      RECT 26.800 -0.500 27.800 0.500 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 9.600 12.500 ;
      RECT 21.600 4.300 30.400 5.300 ;
      RECT 0.800 6.700 22.600 7.700 ;
      RECT 29.400 4.300 30.400 10.100 ;
      RECT 6.000 6.700 22.600 10.100 ;
      RECT 0.800 11.500 12.200 12.500 ;
      RECT 16.400 6.700 22.600 19.700 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 11.200 13.900 22.600 17.300 ;
      RECT 26.800 13.900 27.800 19.700 ;
      RECT 26.800 16.300 30.400 19.700 ;
      RECT 0.800 18.700 1.800 22.100 ;
      RECT 6.000 18.700 7.000 24.500 ;
      RECT 16.400 18.700 30.400 19.700 ;
      RECT 0.800 21.100 7.000 22.100 ;
      RECT 11.200 21.100 14.800 24.500 ;
      RECT 21.600 18.700 25.200 22.100 ;
      RECT 6.000 23.500 14.800 24.500 ;
      RECT 24.200 18.700 25.200 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END LTGG

MACRO LTPFF
  CLASS CORE ;
  FOREIGN LTPFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 36.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 13.900 22.600 14.900 ; # D|0.0@0
    END
  END D
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 6.700 35.600 10.100 ; # PN|0.0@0
    END
  END PN
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 11.500 27.800 12.500 ; # S|0.0@0
    END
  END S
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # QN|0.0@0
      RECT 6.000 13.900 7.000 19.700 ; # QN|0.0@1
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 36.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 36.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 12.200 12.500 ;
      RECT 26.800 6.700 33.000 7.700 ;
      RECT 6.000 9.100 25.200 12.500 ;
      RECT 29.400 6.700 33.000 22.100 ;
      RECT 8.600 9.100 20.000 14.900 ;
      RECT 24.200 13.900 35.600 22.100 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 13.800 9.100 20.000 22.100 ;
      RECT 8.600 18.700 35.600 19.700 ;
      RECT 11.200 18.700 35.600 22.100 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 14.800 0.500 ;
      RECT 34.600 -0.500 35.600 0.500 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 11.200 4.300 14.800 5.300 ;
      RECT 21.600 4.300 35.600 5.300 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 16.400 6.700 33.000 7.700 ;
      RECT 0.800 9.100 27.800 10.100 ;
      RECT 32.000 9.100 35.600 10.100 ;
      RECT 6.000 9.100 25.200 12.500 ;
      RECT 29.400 11.500 33.000 14.900 ;
      RECT 3.400 13.900 7.000 14.900 ;
      RECT 11.200 9.100 20.000 14.900 ;
      RECT 24.200 13.900 35.600 14.900 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 13.800 9.100 20.000 24.500 ;
      RECT 24.200 13.900 27.800 24.500 ;
      RECT 32.000 13.900 35.600 24.500 ;
      RECT 6.000 18.700 35.600 19.700 ;
      RECT 6.000 6.700 7.000 22.100 ;
      RECT 11.200 18.700 35.600 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 13.800 18.700 35.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
  END
END LTPFF

MACRO LTQTFF
  CLASS CORE ;
  FOREIGN LTQTFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 41.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 9.100 40.800 12.500 ; # OE|0.0@0
    END
  END OE
  PIN L
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # L|0.0@0
    END
  END L
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 9.100 25.200 14.900 ; # Q|0.0@0
    END
  END Q
  PIN QT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 9.100 35.600 10.100 ; # QT|0.0@0
    END
  END QT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 41.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 41.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 25.200 7.700 ;
      RECT 29.400 6.700 40.800 7.700 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 11.200 6.700 20.000 22.100 ;
      RECT 29.400 6.700 33.000 19.700 ;
      RECT 37.200 6.700 38.200 19.700 ;
      RECT 3.400 11.500 20.000 12.500 ;
      RECT 29.400 11.500 38.200 19.700 ;
      RECT 11.200 13.900 22.600 17.300 ;
      RECT 11.200 16.300 25.200 17.300 ;
      RECT 3.400 18.700 20.000 19.700 ;
      RECT 24.200 18.700 38.200 19.700 ;
      RECT 8.600 18.700 20.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 26.800 -0.500 27.800 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 19.000 4.300 27.800 7.700 ;
      RECT 37.200 4.300 40.800 7.700 ;
      RECT 3.400 6.700 40.800 7.700 ;
      RECT 0.800 9.100 22.600 10.100 ;
      RECT 26.800 6.700 33.000 22.100 ;
      RECT 37.200 4.300 38.200 22.100 ;
      RECT 0.800 9.100 17.400 12.500 ;
      RECT 26.800 11.500 40.800 12.500 ;
      RECT 3.400 4.300 7.000 24.500 ;
      RECT 11.200 4.300 14.800 22.100 ;
      RECT 21.600 13.900 22.600 17.300 ;
      RECT 26.800 11.500 38.200 22.100 ;
      RECT 11.200 16.300 17.400 22.100 ;
      RECT 21.600 16.300 38.200 17.300 ;
      RECT 3.400 18.700 20.000 22.100 ;
      RECT 24.200 16.300 38.200 22.100 ;
      RECT 0.800 23.500 12.200 24.500 ;
      RECT 16.400 18.700 20.000 24.500 ;
      RECT 26.800 4.300 27.800 24.500 ;
      RECT 39.800 23.500 40.800 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 16.400 28.300 20.000 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
  END
END LTQTFF

MACRO LTQTGG
  CLASS CORE ;
  FOREIGN LTQTGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 49.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # D|0.0@0
    END
  END D
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 9.100 48.600 12.500 ; # OE|0.0@0
    END
  END OE
  PIN L
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # L|0.0@0
    END
  END L
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 27.800 7.700 ; # Q|0.0@0
      RECT 26.800 6.700 27.800 14.900 ; # Q|0.0@1
      RECT 26.800 13.900 30.400 14.900 ; # Q|0.0@2
      RECT 29.400 13.900 30.400 19.700 ; # Q|0.0@3
    END
  END Q
  PIN QT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.200 11.500 38.200 14.900 ; # QT|0.0@0
    END
  END QT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 49.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 49.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 22.600 10.100 ;
      RECT 29.400 6.700 46.000 10.100 ;
      RECT 3.400 9.100 25.200 10.100 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 11.200 9.100 25.200 19.700 ;
      RECT 32.000 6.700 33.000 22.100 ;
      RECT 39.800 6.700 46.000 17.300 ;
      RECT 3.400 16.300 25.200 19.700 ;
      RECT 37.200 16.300 46.000 17.300 ;
      RECT 32.000 18.700 38.200 22.100 ;
      RECT 42.400 6.700 46.000 22.100 ;
      RECT 8.600 16.300 22.600 22.100 ;
      RECT 29.400 21.100 46.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 47.600 -0.500 48.600 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 19.000 4.300 48.600 5.300 ;
      RECT 3.400 4.300 7.000 22.100 ;
      RECT 11.200 6.700 22.600 22.100 ;
      RECT 29.400 4.300 46.000 7.700 ;
      RECT 3.400 9.100 25.200 10.100 ;
      RECT 29.400 4.300 43.400 10.100 ;
      RECT 47.600 9.100 48.600 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 9.100 25.200 14.900 ;
      RECT 29.400 4.300 35.600 12.500 ;
      RECT 39.800 11.500 46.000 24.500 ;
      RECT 32.000 4.300 35.600 22.100 ;
      RECT 3.400 16.300 22.600 22.100 ;
      RECT 26.800 16.300 48.600 17.300 ;
      RECT 3.400 18.700 25.200 22.100 ;
      RECT 29.400 16.300 48.600 19.700 ;
      RECT 29.400 16.300 46.000 22.100 ;
      RECT 8.600 16.300 9.600 24.500 ;
      RECT 13.800 4.300 14.800 24.500 ;
      RECT 24.200 18.700 25.200 24.500 ;
      RECT 34.600 16.300 46.000 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 45.000 28.300 48.600 29.300 ;
  END
END LTQTGG

MACRO LTZFF
  CLASS CORE ;
  FOREIGN LTZFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 36.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN S
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # S|0.0@0
    END
  END S
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 16.300 25.200 17.300 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 6.700 35.600 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 36.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 36.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 11.200 6.700 33.000 14.900 ;
      RECT 3.400 9.100 33.000 12.500 ;
      RECT 3.400 16.300 22.600 19.700 ;
      RECT 29.400 6.700 33.000 22.100 ;
      RECT 3.400 18.700 25.200 19.700 ;
      RECT 3.400 16.300 9.600 22.100 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 24.200 21.100 35.600 22.100 ;
    LAYER cont2 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 19.000 4.300 20.000 5.300 ;
      RECT 24.200 4.300 25.200 14.900 ;
      RECT 29.400 4.300 30.400 24.500 ;
      RECT 3.400 4.300 7.000 24.500 ;
      RECT 11.200 4.300 14.800 19.700 ;
      RECT 24.200 6.700 35.600 10.100 ;
      RECT 11.200 9.100 35.600 10.100 ;
      RECT 0.800 11.500 20.000 12.500 ;
      RECT 24.200 6.700 33.000 14.900 ;
      RECT 11.200 13.900 33.000 14.900 ;
      RECT 3.400 16.300 22.600 19.700 ;
      RECT 29.400 6.700 33.000 24.500 ;
      RECT 3.400 18.700 33.000 19.700 ;
      RECT 3.400 16.300 9.600 24.500 ;
      RECT 16.400 9.100 20.000 22.100 ;
      RECT 24.200 21.100 35.600 24.500 ;
      RECT 0.800 23.500 9.600 24.500 ;
      RECT 21.600 23.500 35.600 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END LTZFF

MACRO MUX2DD
  CLASS CORE ;
  FOREIGN MUX2DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 6.700 22.600 7.700 ; # Q|0.0@0
      RECT 19.000 6.700 20.000 14.900 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 14.800 10.100 ;
      RECT 3.400 9.100 17.400 10.100 ;
      RECT 3.400 9.100 9.600 17.300 ;
      RECT 13.800 9.100 17.400 12.500 ;
      RECT 16.400 9.100 17.400 22.100 ;
      RECT 0.800 16.300 22.600 17.300 ;
      RECT 0.800 16.300 4.400 19.700 ;
      RECT 8.600 16.300 22.600 19.700 ;
      RECT 8.600 6.700 9.600 22.100 ;
      RECT 13.800 16.300 17.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 22.600 5.300 ;
      RECT 8.600 4.300 14.800 10.100 ;
      RECT 21.600 4.300 22.600 12.500 ;
      RECT 3.400 9.100 17.400 10.100 ;
      RECT 0.800 11.500 9.600 12.500 ;
      RECT 13.800 9.100 17.400 12.500 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 9.100 17.400 24.500 ;
      RECT 0.800 16.300 22.600 19.700 ;
      RECT 6.000 16.300 17.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 16.300 17.400 24.500 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END MUX2DD

MACRO MUX2FF
  CLASS CORE ;
  FOREIGN MUX2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 10.100 ; # Q|0.0@0
      RECT 21.600 9.100 25.200 10.100 ; # Q|0.0@1
      RECT 21.600 9.100 22.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 22.600 7.700 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 6.700 20.000 14.900 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 6.700 17.400 17.300 ;
      RECT 6.000 16.300 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 20.000 7.700 ;
      RECT 24.200 4.300 25.200 12.500 ;
      RECT 6.000 6.700 25.200 7.700 ;
      RECT 0.800 9.100 4.400 12.500 ;
      RECT 8.600 4.300 12.200 12.500 ;
      RECT 16.400 4.300 20.000 14.900 ;
      RECT 8.600 11.500 20.000 12.500 ;
      RECT 3.400 9.100 4.400 19.700 ;
      RECT 8.600 4.300 9.600 24.500 ;
      RECT 8.600 16.300 12.200 22.100 ;
      RECT 16.400 4.300 17.400 17.300 ;
      RECT 21.600 16.300 22.600 19.700 ;
      RECT 6.000 21.100 12.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 21.100 9.600 24.500 ;
      RECT 13.800 23.500 20.000 24.500 ;
      RECT 24.200 23.500 25.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END MUX2FF

MACRO MUX2GG
  CLASS CORE ;
  FOREIGN MUX2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 11.500 27.800 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 9.100 25.200 19.700 ; # Q|0.0@0
      RECT 21.600 16.300 25.200 17.300 ; # Q|0.0@1
      RECT 19.000 18.700 20.000 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 20.000 12.500 ;
      RECT 24.200 6.700 25.200 7.700 ;
      RECT 3.400 9.100 20.000 12.500 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 6.700 20.000 17.300 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 6.700 17.400 19.700 ;
      RECT 6.000 6.700 9.600 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 20.000 5.300 ;
      RECT 26.800 4.300 27.800 5.300 ;
      RECT 6.000 4.300 17.400 12.500 ;
      RECT 21.600 6.700 25.200 10.100 ;
      RECT 0.800 9.100 25.200 10.100 ;
      RECT 0.800 9.100 22.600 12.500 ;
      RECT 26.800 11.500 27.800 12.500 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 9.100 22.600 14.900 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 9.100 20.000 19.700 ;
      RECT 24.200 16.300 25.200 22.100 ;
      RECT 16.400 18.700 25.200 19.700 ;
      RECT 6.000 4.300 9.600 22.100 ;
      RECT 19.000 9.100 20.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END MUX2GG

MACRO MUX2HH
  CLASS CORE ;
  FOREIGN MUX2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 10.100 ; # Q|0.0@0
      RECT 24.200 9.100 27.800 10.100 ; # Q|0.0@1
      RECT 26.800 9.100 27.800 17.300 ; # Q|0.0@2
      RECT 21.600 16.300 22.600 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 26.800 6.700 27.800 7.700 ;
      RECT 3.400 6.700 9.600 22.100 ;
      RECT 29.400 11.500 30.400 22.100 ;
      RECT 3.400 16.300 20.000 22.100 ;
      RECT 3.400 18.700 30.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 14.800 5.300 ;
      RECT 24.200 4.300 25.200 12.500 ;
      RECT 29.400 4.300 30.400 5.300 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 16.400 6.700 20.000 14.900 ;
      RECT 24.200 6.700 27.800 7.700 ;
      RECT 3.400 6.700 9.600 22.100 ;
      RECT 0.800 11.500 25.200 12.500 ;
      RECT 29.400 11.500 30.400 14.900 ;
      RECT 16.400 11.500 22.600 14.900 ;
      RECT 0.800 16.300 17.400 22.100 ;
      RECT 21.600 11.500 22.600 24.500 ;
      RECT 26.800 16.300 27.800 24.500 ;
      RECT 0.800 18.700 27.800 19.700 ;
      RECT 21.600 18.700 27.800 24.500 ;
      RECT 0.800 16.300 1.800 24.500 ;
      RECT 11.200 16.300 12.200 24.500 ;
      RECT 19.000 23.500 30.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
  END
END MUX2HH

MACRO MUX2NEDD
  CLASS CORE ;
  FOREIGN MUX2NEDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 20.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 6.700 20.000 22.100 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 20.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 20.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 11.200 6.700 17.400 10.100 ;
      RECT 3.400 11.500 12.200 12.500 ;
      RECT 16.400 6.700 17.400 22.100 ;
      RECT 11.200 13.900 17.400 22.100 ;
      RECT 3.400 16.300 17.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 9.600 7.700 ;
      RECT 19.000 4.300 20.000 7.700 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 0.800 11.500 12.200 12.500 ;
      RECT 16.400 6.700 17.400 24.500 ;
      RECT 3.400 4.300 7.000 22.100 ;
      RECT 11.200 13.900 17.400 24.500 ;
      RECT 3.400 16.300 17.400 22.100 ;
      RECT 3.400 21.100 20.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 21.100 20.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 17.400 29.300 ;
  END
END MUX2NEDD

MACRO MUX2NEFF
  CLASS CORE ;
  FOREIGN MUX2NEFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 6.700 22.600 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 20.000 7.700 ;
      RECT 3.400 9.100 9.600 17.300 ;
      RECT 13.800 6.700 20.000 12.500 ;
      RECT 3.400 11.500 20.000 12.500 ;
      RECT 16.400 6.700 20.000 14.900 ;
      RECT 3.400 16.300 12.200 17.300 ;
      RECT 16.400 6.700 17.400 17.300 ;
      RECT 6.000 16.300 12.200 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 22.600 10.100 ;
      RECT 3.400 9.100 22.600 10.100 ;
      RECT 0.800 11.500 20.000 12.500 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 4.300 20.000 14.900 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 4.300 17.400 17.300 ;
      RECT 21.600 16.300 22.600 19.700 ;
      RECT 6.000 16.300 12.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END MUX2NEFF

MACRO MUX2NEGG
  CLASS CORE ;
  FOREIGN MUX2NEGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 6.700 22.600 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 20.000 7.700 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 13.800 6.700 20.000 12.500 ;
      RECT 3.400 11.500 20.000 12.500 ;
      RECT 16.400 6.700 20.000 14.900 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 6.700 17.400 17.300 ;
      RECT 6.000 16.300 12.200 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 19.000 -0.500 25.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 22.600 10.100 ;
      RECT 3.400 9.100 22.600 10.100 ;
      RECT 0.800 11.500 20.000 12.500 ;
      RECT 3.400 9.100 9.600 19.700 ;
      RECT 16.400 4.300 20.000 17.300 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 16.300 22.600 17.300 ;
      RECT 19.000 16.300 22.600 19.700 ;
      RECT 6.000 16.300 12.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END MUX2NEGG

MACRO MUX2NEHH
  CLASS CORE ;
  FOREIGN MUX2NEHH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 10.100 ; # Y1|0.0@0
    END
  END Y1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 16.400 6.700 22.600 19.700 ;
      RECT 3.400 6.700 9.600 19.700 ;
      RECT 3.400 11.500 12.200 19.700 ;
      RECT 3.400 18.700 22.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 14.800 0.500 ;
      RECT 19.000 -0.500 25.200 0.500 ;
      RECT 0.800 4.300 12.200 7.700 ;
      RECT 16.400 4.300 25.200 5.300 ;
      RECT 16.400 4.300 22.600 19.700 ;
      RECT 3.400 4.300 9.600 19.700 ;
      RECT 13.800 9.100 22.600 12.500 ;
      RECT 0.800 11.500 22.600 12.500 ;
      RECT 3.400 11.500 12.200 19.700 ;
      RECT 3.400 18.700 22.600 19.700 ;
      RECT 21.600 21.100 25.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 24.200 21.100 25.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END MUX2NEHH

MACRO MUX4DD
  CLASS CORE ;
  FOREIGN MUX4DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 67.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 11.500 17.400 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 11.500 33.000 12.500 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 11.500 35.600 14.900 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 45.000 11.500 46.000 12.500 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 13.900 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@0
    END
  END B
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 13.900 56.400 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 65.800 6.700 66.800 19.700 ; # Q|0.0@0
      RECT 60.600 16.300 61.600 17.300 ; # Q|0.0@1
      RECT 55.400 18.700 59.000 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 67.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 67.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 6.000 6.700 64.200 7.700 ;
      RECT 0.800 9.100 46.000 10.100 ;
      RECT 50.200 6.700 64.200 12.500 ;
      RECT 3.400 9.100 7.000 19.700 ;
      RECT 11.200 6.700 14.800 17.300 ;
      RECT 19.000 6.700 30.400 12.500 ;
      RECT 42.400 6.700 43.400 22.100 ;
      RECT 3.400 13.900 14.800 17.300 ;
      RECT 21.600 13.900 33.000 22.100 ;
      RECT 42.400 13.900 53.800 22.100 ;
      RECT 58.000 6.700 64.200 14.900 ;
      RECT 0.800 16.300 53.800 17.300 ;
      RECT 63.200 6.700 64.200 22.100 ;
      RECT 0.800 16.300 9.600 19.700 ;
      RECT 13.800 16.300 53.800 22.100 ;
      RECT 60.600 18.700 64.200 22.100 ;
      RECT 6.000 21.100 66.800 22.100 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 20.000 0.500 ;
      RECT 32.000 -0.500 35.600 0.500 ;
      RECT 39.800 -0.500 46.000 0.500 ;
      RECT 55.400 -0.500 56.400 0.500 ;
      RECT 0.800 4.300 66.800 5.300 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 6.000 4.300 66.800 7.700 ;
      RECT 6.000 4.300 9.600 10.100 ;
      RECT 13.800 4.300 30.400 10.100 ;
      RECT 39.800 4.300 66.800 10.100 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 11.200 11.500 12.200 17.300 ;
      RECT 19.000 4.300 30.400 12.500 ;
      RECT 39.800 4.300 43.400 24.500 ;
      RECT 47.600 4.300 48.600 24.500 ;
      RECT 52.800 4.300 64.200 12.500 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 21.600 13.900 35.600 19.700 ;
      RECT 39.800 13.900 51.200 24.500 ;
      RECT 58.000 4.300 64.200 14.900 ;
      RECT 0.800 16.300 4.400 19.700 ;
      RECT 8.600 13.900 12.200 17.300 ;
      RECT 16.400 16.300 51.200 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 13.800 18.700 56.400 19.700 ;
      RECT 60.600 18.700 61.600 24.500 ;
      RECT 65.800 18.700 66.800 22.100 ;
      RECT 6.000 21.100 27.800 24.500 ;
      RECT 32.000 21.100 61.600 24.500 ;
      RECT 6.000 23.500 64.200 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
      RECT 63.200 28.300 64.200 29.300 ;
  END
END MUX4DD

MACRO MUX4FF
  CLASS CORE ;
  FOREIGN MUX4FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 78.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 9.100 20.000 10.100 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 13.900 30.400 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 9.100 40.800 10.100 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 11.500 48.600 14.900 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 9.100 53.800 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 76.200 6.700 77.200 22.100 ; # Q|0.0@0
      RECT 60.600 21.100 61.600 22.100 ; # Q|0.0@1
      RECT 65.800 21.100 66.800 22.100 ; # Q|0.0@2
      RECT 71.000 21.100 77.200 22.100 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 78.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 78.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 38.200 7.700 ;
      RECT 42.400 6.700 59.000 7.700 ;
      RECT 63.200 6.700 74.600 14.900 ;
      RECT 0.800 9.100 1.800 19.700 ;
      RECT 6.000 6.700 9.600 22.100 ;
      RECT 13.800 6.700 17.400 19.700 ;
      RECT 21.600 6.700 30.400 12.500 ;
      RECT 34.600 6.700 38.200 14.900 ;
      RECT 42.400 6.700 46.000 22.100 ;
      RECT 58.000 9.100 74.600 14.900 ;
      RECT 0.800 11.500 9.600 17.300 ;
      RECT 13.800 11.500 30.400 12.500 ;
      RECT 34.600 11.500 46.000 14.900 ;
      RECT 0.800 13.900 17.400 17.300 ;
      RECT 24.200 6.700 27.800 22.100 ;
      RECT 55.400 13.900 74.600 14.900 ;
      RECT 0.800 16.300 33.000 17.300 ;
      RECT 37.200 16.300 59.000 22.100 ;
      RECT 63.200 6.700 64.200 22.100 ;
      RECT 68.400 6.700 74.600 19.700 ;
      RECT 13.800 16.300 20.000 19.700 ;
      RECT 24.200 18.700 74.600 19.700 ;
      RECT 6.000 21.100 14.800 22.100 ;
      RECT 24.200 18.700 59.000 22.100 ;
      RECT 68.400 6.700 69.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 34.600 -0.500 35.600 0.500 ;
      RECT 52.800 -0.500 53.800 0.500 ;
      RECT 76.200 -0.500 77.200 0.500 ;
      RECT 6.000 4.300 38.200 7.700 ;
      RECT 42.400 4.300 59.000 5.300 ;
      RECT 63.200 4.300 77.200 5.300 ;
      RECT 42.400 4.300 56.400 7.700 ;
      RECT 63.200 4.300 74.600 7.700 ;
      RECT 0.800 9.100 1.800 19.700 ;
      RECT 6.000 4.300 12.200 10.100 ;
      RECT 21.600 4.300 30.400 10.100 ;
      RECT 34.600 4.300 38.200 17.300 ;
      RECT 45.000 4.300 46.000 24.500 ;
      RECT 58.000 9.100 72.000 14.900 ;
      RECT 0.800 11.500 9.600 17.300 ;
      RECT 13.800 11.500 14.800 19.700 ;
      RECT 19.000 11.500 22.600 12.500 ;
      RECT 29.400 4.300 30.400 12.500 ;
      RECT 34.600 11.500 46.000 14.900 ;
      RECT 58.000 11.500 74.600 14.900 ;
      RECT 0.800 13.900 17.400 17.300 ;
      RECT 34.600 13.900 48.600 14.900 ;
      RECT 52.800 13.900 77.200 14.900 ;
      RECT 0.800 16.300 27.800 17.300 ;
      RECT 32.000 16.300 38.200 17.300 ;
      RECT 42.400 16.300 66.800 19.700 ;
      RECT 71.000 13.900 77.200 19.700 ;
      RECT 6.000 16.300 20.000 19.700 ;
      RECT 24.200 18.700 33.000 22.100 ;
      RECT 37.200 18.700 77.200 19.700 ;
      RECT 6.000 13.900 12.200 24.500 ;
      RECT 24.200 21.100 59.000 22.100 ;
      RECT 63.200 4.300 64.200 22.100 ;
      RECT 68.400 18.700 69.400 22.100 ;
      RECT 76.200 13.900 77.200 22.100 ;
      RECT 3.400 23.500 14.800 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 29.400 21.100 56.400 24.500 ;
      RECT 60.600 23.500 61.600 24.500 ;
      RECT 65.800 23.500 66.800 24.500 ;
      RECT 71.000 23.500 74.600 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 11.200 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
      RECT 45.000 28.300 48.600 29.300 ;
      RECT 55.400 28.300 56.400 29.300 ;
      RECT 60.600 28.300 61.600 29.300 ;
      RECT 65.800 28.300 66.800 29.300 ;
      RECT 71.000 28.300 74.600 29.300 ;
  END
END MUX4FF

MACRO MUX4GG
  CLASS CORE ;
  FOREIGN MUX4GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 85.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 13.900 33.000 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 11.500 43.400 12.500 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 50.200 13.900 51.200 14.900 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 84.000 6.700 85.000 17.300 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 73.600 9.100 82.400 10.100 ; # Q|0.0@0
      RECT 81.400 9.100 82.400 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 85.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 85.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 22.100 ;
      RECT 6.000 6.700 9.600 22.100 ;
      RECT 16.400 6.700 40.800 7.700 ;
      RECT 45.000 6.700 82.400 7.700 ;
      RECT 13.800 9.100 20.000 19.700 ;
      RECT 26.800 6.700 40.800 12.500 ;
      RECT 45.000 6.700 61.600 12.500 ;
      RECT 65.800 6.700 72.000 22.100 ;
      RECT 0.800 11.500 9.600 14.900 ;
      RECT 45.000 11.500 77.200 12.500 ;
      RECT 0.800 13.900 20.000 14.900 ;
      RECT 26.800 6.700 30.400 22.100 ;
      RECT 34.600 6.700 38.200 22.100 ;
      RECT 45.000 6.700 48.600 22.100 ;
      RECT 52.800 13.900 79.800 22.100 ;
      RECT 6.000 16.300 79.800 19.700 ;
      RECT 6.000 18.700 85.000 19.700 ;
      RECT 6.000 13.900 17.400 22.100 ;
      RECT 24.200 18.700 82.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 19.000 -0.500 22.600 0.500 ;
      RECT 37.200 -0.500 40.800 0.500 ;
      RECT 55.400 -0.500 56.400 0.500 ;
      RECT 81.400 -0.500 82.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 8.600 4.300 9.600 24.500 ;
      RECT 13.800 4.300 40.800 5.300 ;
      RECT 45.000 4.300 85.000 5.300 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 6.000 6.700 9.600 24.500 ;
      RECT 16.400 4.300 38.200 7.700 ;
      RECT 45.000 4.300 53.800 7.700 ;
      RECT 58.000 4.300 82.400 7.700 ;
      RECT 13.800 9.100 20.000 17.300 ;
      RECT 24.200 4.300 33.000 10.100 ;
      RECT 37.200 9.100 51.200 10.100 ;
      RECT 55.400 9.100 61.600 17.300 ;
      RECT 65.800 4.300 72.000 10.100 ;
      RECT 3.400 11.500 9.600 14.900 ;
      RECT 26.800 11.500 40.800 12.500 ;
      RECT 45.000 4.300 51.200 12.500 ;
      RECT 55.400 11.500 64.200 17.300 ;
      RECT 76.200 11.500 77.200 22.100 ;
      RECT 3.400 13.900 30.400 14.900 ;
      RECT 34.600 13.900 48.600 24.500 ;
      RECT 55.400 13.900 79.800 17.300 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 6.000 16.300 79.800 17.300 ;
      RECT 84.000 16.300 85.000 19.700 ;
      RECT 6.000 13.900 17.400 19.700 ;
      RECT 21.600 13.900 22.600 19.700 ;
      RECT 26.800 16.300 56.400 24.500 ;
      RECT 60.600 18.700 85.000 19.700 ;
      RECT 16.400 4.300 17.400 22.100 ;
      RECT 24.200 21.100 56.400 24.500 ;
      RECT 60.600 18.700 82.400 22.100 ;
      RECT 3.400 23.500 12.200 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 24.200 23.500 59.000 24.500 ;
      RECT 63.200 11.500 64.200 24.500 ;
      RECT 68.400 13.900 69.400 24.500 ;
      RECT 73.600 13.900 74.600 24.500 ;
      RECT 78.800 13.900 79.800 24.500 ;
      RECT 84.000 23.500 85.000 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 37.200 28.300 46.000 29.300 ;
      RECT 52.800 28.300 53.800 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
      RECT 68.400 28.300 69.400 29.300 ;
      RECT 78.800 28.300 79.800 29.300 ;
  END
END MUX4GG

MACRO MUX4HH
  CLASS CORE ;
  FOREIGN MUX4HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 135.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 11.500 30.400 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 11.500 51.200 12.500 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 60.600 11.500 61.600 12.500 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 81.400 11.500 82.400 12.500 ; # Y3|0.0@0
      RECT 86.600 11.500 90.200 12.500 ; # Y3|0.0@1
      RECT 78.800 13.900 79.800 14.900 ; # Y3|0.0@2
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 12.500 ; # B|0.0@0
    END
  END B
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 117.800 11.500 118.800 12.500 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 128.200 6.700 129.200 7.700 ; # Q|0.0@0
      RECT 133.400 6.700 134.400 22.100 ; # Q|0.0@1
      RECT 99.600 21.100 100.600 22.100 ; # Q|0.0@2
      RECT 110.000 21.100 111.000 22.100 ; # Q|0.0@3
      RECT 115.200 21.100 116.200 22.100 ; # Q|0.0@4
      RECT 128.200 21.100 129.200 22.100 ; # Q|0.0@5
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 135.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 135.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 19.000 6.700 59.000 7.700 ;
      RECT 63.200 6.700 126.600 7.700 ;
      RECT 130.800 6.700 131.800 22.100 ;
      RECT 3.400 9.100 4.400 17.300 ;
      RECT 8.600 9.100 12.200 19.700 ;
      RECT 16.400 9.100 22.600 19.700 ;
      RECT 29.400 6.700 33.000 10.100 ;
      RECT 45.000 6.700 48.600 10.100 ;
      RECT 55.400 6.700 59.000 22.100 ;
      RECT 63.200 6.700 72.000 12.500 ;
      RECT 76.200 6.700 85.000 10.100 ;
      RECT 91.800 9.100 131.800 10.100 ;
      RECT 32.000 6.700 33.000 22.100 ;
      RECT 45.000 6.700 46.000 22.100 ;
      RECT 76.200 6.700 79.800 12.500 ;
      RECT 84.000 6.700 85.000 12.500 ;
      RECT 91.800 6.700 116.200 19.700 ;
      RECT 120.400 9.100 131.800 19.700 ;
      RECT 3.400 13.900 22.600 17.300 ;
      RECT 68.400 6.700 72.000 22.100 ;
      RECT 76.200 6.700 77.200 22.100 ;
      RECT 89.200 13.900 131.800 19.700 ;
      RECT 3.400 16.300 72.000 17.300 ;
      RECT 76.200 16.300 131.800 19.700 ;
      RECT 8.600 18.700 131.800 19.700 ;
      RECT 32.000 18.700 98.000 22.100 ;
      RECT 102.200 6.700 108.400 22.100 ;
      RECT 112.600 6.700 113.600 22.100 ;
      RECT 117.800 13.900 126.600 22.100 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 45.000 -0.500 46.000 0.500 ;
      RECT 89.200 -0.500 92.800 0.500 ;
      RECT 117.800 -0.500 118.800 0.500 ;
      RECT 6.000 4.300 7.000 5.300 ;
      RECT 13.800 4.300 14.800 5.300 ;
      RECT 19.000 4.300 59.000 5.300 ;
      RECT 73.600 4.300 77.200 5.300 ;
      RECT 91.800 4.300 92.800 5.300 ;
      RECT 102.200 4.300 134.400 5.300 ;
      RECT 19.000 4.300 20.000 19.700 ;
      RECT 24.200 4.300 59.000 7.700 ;
      RECT 63.200 6.700 69.400 22.100 ;
      RECT 84.000 6.700 85.000 14.900 ;
      RECT 99.600 6.700 126.600 7.700 ;
      RECT 130.800 4.300 131.800 24.500 ;
      RECT 0.800 9.100 4.400 17.300 ;
      RECT 8.600 9.100 12.200 10.100 ;
      RECT 16.400 9.100 22.600 19.700 ;
      RECT 26.800 4.300 33.000 10.100 ;
      RECT 45.000 4.300 51.200 10.100 ;
      RECT 55.400 9.100 72.000 10.100 ;
      RECT 84.000 9.100 87.600 10.100 ;
      RECT 91.800 9.100 95.400 24.500 ;
      RECT 99.600 6.700 121.400 10.100 ;
      RECT 125.600 9.100 131.800 19.700 ;
      RECT 8.600 9.100 9.600 19.700 ;
      RECT 29.400 4.300 33.000 19.700 ;
      RECT 45.000 4.300 48.600 19.700 ;
      RECT 55.400 4.300 59.000 22.100 ;
      RECT 63.200 9.100 72.000 22.100 ;
      RECT 76.200 11.500 79.800 12.500 ;
      RECT 89.200 11.500 116.200 14.900 ;
      RECT 120.400 11.500 131.800 19.700 ;
      RECT 0.800 13.900 9.600 17.300 ;
      RECT 13.800 13.900 72.000 14.900 ;
      RECT 76.200 11.500 77.200 14.900 ;
      RECT 81.400 13.900 131.800 14.900 ;
      RECT 13.800 13.900 48.600 19.700 ;
      RECT 52.800 13.900 72.000 22.100 ;
      RECT 78.800 16.300 82.400 24.500 ;
      RECT 86.600 13.900 87.600 24.500 ;
      RECT 91.800 13.900 131.800 19.700 ;
      RECT 3.400 18.700 72.000 19.700 ;
      RECT 78.800 18.700 131.800 19.700 ;
      RECT 32.000 4.300 33.000 22.100 ;
      RECT 50.200 21.100 98.000 22.100 ;
      RECT 102.200 4.300 108.400 24.500 ;
      RECT 112.600 4.300 113.600 24.500 ;
      RECT 117.800 13.900 126.600 24.500 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 9.600 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 24.200 23.500 25.200 24.500 ;
      RECT 29.400 23.500 30.400 24.500 ;
      RECT 34.600 23.500 35.600 24.500 ;
      RECT 39.800 23.500 40.800 24.500 ;
      RECT 45.000 23.500 46.000 24.500 ;
      RECT 50.200 18.700 53.800 24.500 ;
      RECT 58.000 4.300 59.000 24.500 ;
      RECT 63.200 6.700 64.200 24.500 ;
      RECT 68.400 6.700 69.400 24.500 ;
      RECT 73.600 23.500 134.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 9.600 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
      RECT 63.200 28.300 64.200 29.300 ;
      RECT 68.400 28.300 69.400 29.300 ;
      RECT 73.600 28.300 77.200 29.300 ;
      RECT 81.400 28.300 82.400 29.300 ;
      RECT 86.600 28.300 87.600 29.300 ;
      RECT 94.400 28.300 95.400 29.300 ;
      RECT 104.800 28.300 105.800 29.300 ;
      RECT 115.200 28.300 118.800 29.300 ;
      RECT 128.200 28.300 129.200 29.300 ;
  END
END MUX4HH

MACRO MUX4NEDD
  CLASS CORE ;
  FOREIGN MUX4NEDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 65.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 13.900 30.400 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 11.500 43.400 14.900 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 45.000 11.500 46.000 14.900 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 10.100 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 63.200 6.700 64.200 19.700 ; # Q|0.0@0
      RECT 58.000 18.700 64.200 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 65.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 65.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ;
      RECT 8.600 6.700 59.000 7.700 ;
      RECT 6.000 9.100 12.200 17.300 ;
      RECT 16.400 6.700 38.200 10.100 ;
      RECT 50.200 6.700 59.000 17.300 ;
      RECT 0.800 11.500 22.600 14.900 ;
      RECT 26.800 6.700 38.200 12.500 ;
      RECT 50.200 11.500 61.600 17.300 ;
      RECT 0.800 13.900 27.800 14.900 ;
      RECT 32.000 6.700 38.200 14.900 ;
      RECT 6.000 11.500 22.600 17.300 ;
      RECT 26.800 16.300 33.000 22.100 ;
      RECT 37.200 16.300 61.600 17.300 ;
      RECT 6.000 9.100 9.600 22.100 ;
      RECT 19.000 18.700 56.400 19.700 ;
      RECT 6.000 21.100 46.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 12.200 0.500 ;
      RECT 52.800 -0.500 53.800 0.500 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 8.600 4.300 38.200 7.700 ;
      RECT 42.400 4.300 46.000 7.700 ;
      RECT 52.800 4.300 53.800 19.700 ;
      RECT 63.200 4.300 64.200 7.700 ;
      RECT 0.800 4.300 1.800 19.700 ;
      RECT 6.000 6.700 59.000 7.700 ;
      RECT 6.000 6.700 12.200 22.100 ;
      RECT 16.400 6.700 43.400 10.100 ;
      RECT 50.200 6.700 59.000 17.300 ;
      RECT 0.800 11.500 22.600 17.300 ;
      RECT 26.800 4.300 38.200 12.500 ;
      RECT 50.200 11.500 61.600 17.300 ;
      RECT 0.800 13.900 27.800 17.300 ;
      RECT 32.000 13.900 61.600 17.300 ;
      RECT 0.800 16.300 61.600 17.300 ;
      RECT 6.000 16.300 56.400 19.700 ;
      RECT 60.600 11.500 61.600 19.700 ;
      RECT 6.000 16.300 46.000 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 11.500 17.400 24.500 ;
      RECT 21.600 16.300 30.400 24.500 ;
      RECT 34.600 4.300 35.600 24.500 ;
      RECT 39.800 23.500 48.600 24.500 ;
      RECT 52.800 23.500 53.800 24.500 ;
      RECT 58.000 23.500 59.000 24.500 ;
      RECT 63.200 23.500 64.200 24.500 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
      RECT 63.200 28.300 64.200 29.300 ;
  END
END MUX4NEDD

MACRO MUX4NEFF
  CLASS CORE ;
  FOREIGN MUX4NEFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 72.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 11.500 30.400 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 11.500 43.400 12.500 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 11.500 48.600 12.500 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 63.200 9.100 69.400 10.100 ; # Q|0.0@0
      RECT 68.400 9.100 69.400 14.900 ; # Q|0.0@1
      RECT 65.800 18.700 66.800 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 72.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 72.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 38.200 7.700 ;
      RECT 42.400 6.700 61.600 10.100 ;
      RECT 0.800 6.700 17.400 10.100 ;
      RECT 24.200 6.700 38.200 10.100 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 11.200 6.700 14.800 17.300 ;
      RECT 24.200 6.700 27.800 22.100 ;
      RECT 34.600 6.700 38.200 12.500 ;
      RECT 45.000 6.700 46.000 22.100 ;
      RECT 50.200 6.700 61.600 19.700 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 45.000 13.900 66.800 17.300 ;
      RECT 71.000 13.900 72.000 22.100 ;
      RECT 0.800 16.300 14.800 17.300 ;
      RECT 19.000 16.300 72.000 17.300 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 16.300 9.600 22.100 ;
      RECT 13.800 6.700 14.800 22.100 ;
      RECT 19.000 16.300 64.200 19.700 ;
      RECT 68.400 16.300 72.000 22.100 ;
      RECT 6.000 21.100 46.000 22.100 ;
      RECT 55.400 21.100 72.000 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 26.800 -0.500 27.800 0.500 ;
      RECT 34.600 -0.500 38.200 0.500 ;
      RECT 52.800 -0.500 53.800 0.500 ;
      RECT 71.000 -0.500 72.000 0.500 ;
      RECT 0.800 4.300 38.200 7.700 ;
      RECT 42.400 4.300 61.600 10.100 ;
      RECT 42.400 6.700 69.400 7.700 ;
      RECT 0.800 4.300 17.400 10.100 ;
      RECT 21.600 9.100 64.200 10.100 ;
      RECT 3.400 4.300 7.000 17.300 ;
      RECT 11.200 4.300 17.400 22.100 ;
      RECT 24.200 4.300 38.200 12.500 ;
      RECT 42.400 4.300 46.000 22.100 ;
      RECT 50.200 11.500 66.800 17.300 ;
      RECT 71.000 11.500 72.000 24.500 ;
      RECT 21.600 13.900 27.800 24.500 ;
      RECT 34.600 4.300 35.600 24.500 ;
      RECT 39.800 13.900 66.800 17.300 ;
      RECT 0.800 16.300 72.000 17.300 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 6.000 16.300 64.200 19.700 ;
      RECT 68.400 16.300 72.000 24.500 ;
      RECT 6.000 16.300 48.600 22.100 ;
      RECT 52.800 21.100 72.000 24.500 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 11.200 4.300 12.200 24.500 ;
      RECT 16.400 4.300 17.400 24.500 ;
      RECT 21.600 16.300 38.200 24.500 ;
      RECT 45.000 4.300 46.000 24.500 ;
      RECT 50.200 23.500 72.000 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 34.600 28.300 43.400 29.300 ;
      RECT 50.200 28.300 53.800 29.300 ;
      RECT 60.600 28.300 61.600 29.300 ;
      RECT 65.800 28.300 66.800 29.300 ;
      RECT 71.000 28.300 72.000 29.300 ;
  END
END MUX4NEFF

MACRO MUX4NEGG
  CLASS CORE ;
  FOREIGN MUX4NEGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 80.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 11.500 35.600 12.500 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 11.500 46.000 12.500 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 11.500 53.800 12.500 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 65.800 9.100 72.000 10.100 ; # Q|0.0@0
      RECT 71.000 9.100 72.000 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 80.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 80.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 16.400 6.700 40.800 7.700 ;
      RECT 45.000 6.700 74.600 7.700 ;
      RECT 0.800 9.100 1.800 19.700 ;
      RECT 6.000 9.100 9.600 22.100 ;
      RECT 13.800 9.100 20.000 22.100 ;
      RECT 26.800 6.700 40.800 10.100 ;
      RECT 45.000 6.700 56.400 10.100 ;
      RECT 60.600 6.700 61.600 22.100 ;
      RECT 73.600 6.700 74.600 14.900 ;
      RECT 26.800 6.700 33.000 12.500 ;
      RECT 37.200 6.700 40.800 12.500 ;
      RECT 47.600 6.700 51.200 12.500 ;
      RECT 55.400 6.700 56.400 19.700 ;
      RECT 73.600 11.500 77.200 14.900 ;
      RECT 0.800 13.900 20.000 17.300 ;
      RECT 26.800 6.700 30.400 22.100 ;
      RECT 37.200 6.700 38.200 22.100 ;
      RECT 47.600 6.700 48.600 22.100 ;
      RECT 55.400 13.900 69.400 14.900 ;
      RECT 73.600 13.900 79.800 14.900 ;
      RECT 0.800 16.300 61.600 17.300 ;
      RECT 68.400 13.900 69.400 22.100 ;
      RECT 78.800 13.900 79.800 22.100 ;
      RECT 6.000 16.300 22.600 22.100 ;
      RECT 26.800 18.700 79.800 19.700 ;
      RECT 6.000 21.100 48.600 22.100 ;
      RECT 58.000 18.700 79.800 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 37.200 -0.500 40.800 0.500 ;
      RECT 58.000 -0.500 59.000 0.500 ;
      RECT 78.800 -0.500 79.800 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 8.600 4.300 9.600 5.300 ;
      RECT 13.800 4.300 40.800 5.300 ;
      RECT 45.000 4.300 74.600 7.700 ;
      RECT 78.800 4.300 79.800 5.300 ;
      RECT 16.400 4.300 40.800 7.700 ;
      RECT 0.800 9.100 1.800 19.700 ;
      RECT 6.000 9.100 9.600 22.100 ;
      RECT 13.800 9.100 20.000 22.100 ;
      RECT 24.200 9.100 56.400 10.100 ;
      RECT 60.600 4.300 61.600 22.100 ;
      RECT 65.800 4.300 69.400 22.100 ;
      RECT 73.600 4.300 74.600 24.500 ;
      RECT 26.800 4.300 33.000 24.500 ;
      RECT 37.200 4.300 40.800 12.500 ;
      RECT 45.000 4.300 51.200 19.700 ;
      RECT 55.400 4.300 56.400 19.700 ;
      RECT 60.600 11.500 69.400 22.100 ;
      RECT 73.600 11.500 79.800 22.100 ;
      RECT 0.800 13.900 20.000 17.300 ;
      RECT 24.200 13.900 38.200 24.500 ;
      RECT 42.400 13.900 69.400 19.700 ;
      RECT 0.800 16.300 69.400 17.300 ;
      RECT 6.000 18.700 79.800 19.700 ;
      RECT 6.000 16.300 48.600 22.100 ;
      RECT 58.000 18.700 79.800 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 9.100 9.600 24.500 ;
      RECT 13.800 9.100 14.800 24.500 ;
      RECT 19.000 4.300 20.000 24.500 ;
      RECT 24.200 16.300 40.800 24.500 ;
      RECT 47.600 4.300 48.600 24.500 ;
      RECT 52.800 23.500 53.800 24.500 ;
      RECT 58.000 13.900 59.000 24.500 ;
      RECT 63.200 11.500 64.200 24.500 ;
      RECT 68.400 4.300 69.400 24.500 ;
      RECT 78.800 11.500 79.800 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 37.200 28.300 46.000 29.300 ;
      RECT 52.800 28.300 53.800 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
      RECT 68.400 28.300 69.400 29.300 ;
      RECT 78.800 28.300 79.800 29.300 ;
  END
END MUX4NEGG

MACRO MUX4NEHH
  CLASS CORE ;
  FOREIGN MUX4NEHH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 93.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 12.500 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 11.500 40.800 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 42.400 11.500 43.400 14.900 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 11.500 56.400 12.500 ; # Y3|0.0@0
    END
  END Y3
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 91.800 6.700 92.800 19.700 ; # Q|0.0@0
      RECT 76.200 18.700 77.200 19.700 ; # Q|0.0@1
      RECT 81.400 18.700 82.400 19.700 ; # Q|0.0@2
      RECT 86.600 18.700 87.600 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 93.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 93.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 19.000 6.700 90.200 7.700 ;
      RECT 0.800 9.100 1.800 17.300 ;
      RECT 6.000 9.100 12.200 12.500 ;
      RECT 16.400 9.100 20.000 19.700 ;
      RECT 29.400 6.700 35.600 22.100 ;
      RECT 47.600 6.700 87.600 10.100 ;
      RECT 24.200 11.500 35.600 19.700 ;
      RECT 47.600 6.700 53.800 22.100 ;
      RECT 60.600 11.500 90.200 12.500 ;
      RECT 0.800 13.900 9.600 17.300 ;
      RECT 13.800 13.900 35.600 17.300 ;
      RECT 47.600 13.900 82.400 17.300 ;
      RECT 86.600 11.500 90.200 17.300 ;
      RECT 0.800 16.300 90.200 17.300 ;
      RECT 16.400 16.300 74.600 19.700 ;
      RECT 78.800 6.700 79.800 22.100 ;
      RECT 84.000 16.300 85.000 22.100 ;
      RECT 89.200 11.500 90.200 22.100 ;
      RECT 26.800 16.300 64.200 22.100 ;
      RECT 68.400 6.700 69.400 22.100 ;
      RECT 73.600 6.700 74.600 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 12.200 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 42.400 -0.500 43.400 0.500 ;
      RECT 60.600 -0.500 61.600 0.500 ;
      RECT 81.400 -0.500 82.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 8.600 4.300 12.200 5.300 ;
      RECT 16.400 4.300 92.800 5.300 ;
      RECT 19.000 4.300 92.800 7.700 ;
      RECT 0.800 9.100 1.800 19.700 ;
      RECT 6.000 9.100 12.200 19.700 ;
      RECT 16.400 9.100 35.600 10.100 ;
      RECT 47.600 4.300 87.600 10.100 ;
      RECT 91.800 4.300 92.800 10.100 ;
      RECT 16.400 9.100 20.000 19.700 ;
      RECT 24.200 4.300 35.600 19.700 ;
      RECT 45.000 11.500 53.800 24.500 ;
      RECT 58.000 11.500 90.200 12.500 ;
      RECT 0.800 13.900 82.400 17.300 ;
      RECT 86.600 11.500 90.200 17.300 ;
      RECT 0.800 16.300 90.200 17.300 ;
      RECT 0.800 13.900 74.600 19.700 ;
      RECT 78.800 4.300 79.800 22.100 ;
      RECT 84.000 16.300 85.000 22.100 ;
      RECT 89.200 11.500 90.200 22.100 ;
      RECT 26.800 13.900 74.600 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 26.800 13.900 66.800 24.500 ;
      RECT 71.000 4.300 72.000 24.500 ;
      RECT 76.200 23.500 77.200 24.500 ;
      RECT 81.400 23.500 82.400 24.500 ;
      RECT 86.600 23.500 87.600 24.500 ;
      RECT 91.800 23.500 92.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 34.600 28.300 35.600 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 55.400 28.300 56.400 29.300 ;
      RECT 60.600 28.300 61.600 29.300 ;
      RECT 65.800 28.300 66.800 29.300 ;
      RECT 71.000 28.300 72.000 29.300 ;
      RECT 76.200 28.300 77.200 29.300 ;
      RECT 81.400 28.300 82.400 29.300 ;
      RECT 86.600 28.300 87.600 29.300 ;
      RECT 91.800 28.300 92.800 29.300 ;
  END
END MUX4NEHH

MACRO MUX8GG
  CLASS CORE ;
  FOREIGN MUX8GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 135.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN Y0
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # Y0|0.0@0
    END
  END Y0
  PIN Y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 133.400 11.500 134.400 14.900 ; # Y1|0.0@0
    END
  END Y1
  PIN Y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 11.500 40.800 12.500 ; # Y2|0.0@0
    END
  END Y2
  PIN Y3
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 94.400 9.100 95.400 10.100 ; # Y3|0.0@0
    END
  END Y3
  PIN Y4
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # Y4|0.0@0
    END
  END Y4
  PIN Y5
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 125.600 11.500 126.600 14.900 ; # Y5|0.0@0
    END
  END Y5
  PIN Y6
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 45.000 11.500 46.000 12.500 ; # Y6|0.0@0
    END
  END Y6
  PIN Y7
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 84.000 11.500 85.000 14.900 ; # Y7|0.0@0
    END
  END Y7
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 58.000 6.700 59.000 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 60.600 9.100 61.600 10.100 ; # B|0.0@0
      RECT 60.600 13.900 61.600 14.900 ; # B|0.0@1
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 52.800 11.500 53.800 12.500 ; # C|0.0@0
    END
  END C
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 68.400 9.100 69.400 10.100 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 78.800 9.100 79.800 14.900 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 135.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 135.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 29.400 6.700 56.400 10.100 ;
      RECT 60.600 6.700 111.000 7.700 ;
      RECT 115.200 6.700 118.800 22.100 ;
      RECT 123.000 6.700 129.200 7.700 ;
      RECT 3.400 9.100 7.000 12.500 ;
      RECT 11.200 9.100 56.400 10.100 ;
      RECT 63.200 6.700 66.800 22.100 ;
      RECT 71.000 6.700 77.200 22.100 ;
      RECT 86.600 6.700 92.800 22.100 ;
      RECT 97.000 6.700 111.000 14.900 ;
      RECT 115.200 9.100 124.000 19.700 ;
      RECT 128.200 9.100 131.800 12.500 ;
      RECT 11.200 9.100 38.200 14.900 ;
      RECT 47.600 6.700 51.200 22.100 ;
      RECT 55.400 11.500 77.200 12.500 ;
      RECT 81.400 11.500 82.400 22.100 ;
      RECT 86.600 11.500 124.000 14.900 ;
      RECT 3.400 9.100 4.400 19.700 ;
      RECT 8.600 13.900 59.000 14.900 ;
      RECT 63.200 11.500 77.200 22.100 ;
      RECT 130.800 9.100 131.800 19.700 ;
      RECT 0.800 16.300 25.200 17.300 ;
      RECT 29.400 16.300 105.800 22.100 ;
      RECT 110.000 16.300 126.600 19.700 ;
      RECT 3.400 18.700 131.800 19.700 ;
      RECT 11.200 18.700 121.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 19.000 -0.500 22.600 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 47.600 -0.500 66.800 0.500 ;
      RECT 81.400 -0.500 82.400 0.500 ;
      RECT 91.800 -0.500 98.000 0.500 ;
      RECT 112.600 -0.500 116.200 0.500 ;
      RECT 123.000 -0.500 124.000 0.500 ;
      RECT 128.200 -0.500 129.200 0.500 ;
      RECT 133.400 -0.500 134.400 0.500 ;
      RECT 0.800 4.300 9.600 5.300 ;
      RECT 16.400 4.300 22.600 5.300 ;
      RECT 29.400 4.300 46.000 10.100 ;
      RECT 52.800 4.300 53.800 10.100 ;
      RECT 58.000 4.300 111.000 5.300 ;
      RECT 115.200 4.300 118.800 24.500 ;
      RECT 123.000 4.300 134.400 5.300 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 16.400 4.300 20.000 24.500 ;
      RECT 29.400 6.700 56.400 10.100 ;
      RECT 60.600 4.300 111.000 7.700 ;
      RECT 123.000 4.300 129.200 7.700 ;
      RECT 3.400 9.100 7.000 19.700 ;
      RECT 11.200 9.100 56.400 10.100 ;
      RECT 63.200 4.300 66.800 10.100 ;
      RECT 71.000 4.300 77.200 24.500 ;
      RECT 86.600 4.300 92.800 24.500 ;
      RECT 97.000 4.300 111.000 24.500 ;
      RECT 115.200 9.100 124.000 22.100 ;
      RECT 128.200 9.100 131.800 12.500 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 9.100 38.200 14.900 ;
      RECT 47.600 6.700 51.200 24.500 ;
      RECT 55.400 11.500 61.600 12.500 ;
      RECT 65.800 11.500 77.200 24.500 ;
      RECT 81.400 11.500 82.400 24.500 ;
      RECT 86.600 11.500 124.000 22.100 ;
      RECT 3.400 13.900 59.000 14.900 ;
      RECT 63.200 13.900 77.200 24.500 ;
      RECT 86.600 13.900 126.600 22.100 ;
      RECT 130.800 13.900 134.400 17.300 ;
      RECT 0.800 16.300 25.200 17.300 ;
      RECT 29.400 16.300 126.600 22.100 ;
      RECT 3.400 18.700 131.800 19.700 ;
      RECT 11.200 18.700 131.800 22.100 ;
      RECT 16.400 18.700 118.800 24.500 ;
      RECT 133.400 23.500 134.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
      RECT 37.200 28.300 40.800 29.300 ;
      RECT 45.000 28.300 46.000 29.300 ;
      RECT 50.200 28.300 53.800 29.300 ;
      RECT 58.000 28.300 61.600 29.300 ;
      RECT 65.800 28.300 66.800 29.300 ;
      RECT 71.000 28.300 72.000 29.300 ;
      RECT 76.200 28.300 77.200 29.300 ;
      RECT 86.600 28.300 87.600 29.300 ;
      RECT 97.000 28.300 98.000 29.300 ;
      RECT 102.200 28.300 103.200 29.300 ;
      RECT 110.000 28.300 113.600 29.300 ;
      RECT 123.000 28.300 126.600 29.300 ;
      RECT 133.400 28.300 134.400 29.300 ;
  END
END MUX8GG

MACRO NAND2EE
  CLASS CORE ;
  FOREIGN NAND2EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 7.000 10.100 ; # Q|0.0@0
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END NAND2EE

MACRO NAND2FF
  CLASS CORE ;
  FOREIGN NAND2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 7.000 10.100 ; # Q|0.0@0
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 9.100 7.000 12.500 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 3.400 16.300 4.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END NAND2FF

MACRO NAND2GG
  CLASS CORE ;
  FOREIGN NAND2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 22.100 ; # B|0.0@0
      RECT 11.200 11.500 12.200 22.100 ; # B|0.0@1
      RECT 0.800 21.100 12.200 22.100 ; # B|0.0@2
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@0
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 12.500 ;
    LAYER cont2 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 11.200 4.300 12.200 5.300 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 11.200 11.500 12.200 14.900 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 9.600 29.300 ;
  END
END NAND2GG

MACRO NAND2HH
  CLASS CORE ;
  FOREIGN NAND2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 22.100 ; # B|0.0@0
      RECT 11.200 11.500 12.200 22.100 ; # B|0.0@1
      RECT 0.800 21.100 12.200 22.100 ; # B|0.0@2
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 7.700 ; # Q|0.0@0
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@1
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 11.200 4.300 12.200 5.300 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 11.200 11.500 12.200 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END NAND2HH

MACRO NAND2II
  CLASS CORE ;
  FOREIGN NAND2II 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 19.700 ; # A|0.0@0
      RECT 16.400 13.900 17.400 19.700 ; # A|0.0@1
      RECT 6.000 18.700 17.400 19.700 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 12.500 ; # B|0.0@0
      RECT 11.200 6.700 12.200 12.500 ; # B|0.0@1
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 10.100 ; # Q|0.0@0
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@1
      RECT 8.600 9.100 9.600 14.900 ; # Q|0.0@2
      RECT 13.800 9.100 17.400 10.100 ; # Q|0.0@3
      RECT 13.800 9.100 14.800 14.900 ; # Q|0.0@4
      RECT 11.200 16.300 12.200 17.300 ; # Q|0.0@5
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 5.700 21.600 7.300 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 16.400 11.500 17.400 12.500 ;
      RECT 11.200 13.900 12.200 14.900 ;
      RECT 8.600 16.300 9.600 17.300 ;
      RECT 13.800 16.300 14.800 17.300 ;
      RECT 6.000 21.100 7.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 11.200 4.300 12.200 5.300 ;
      RECT 16.400 4.300 17.400 14.900 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 13.800 6.700 17.400 7.700 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 11.200 13.900 12.200 14.900 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 8.600 16.300 9.600 17.300 ;
      RECT 13.800 16.300 14.800 17.300 ;
      RECT 6.000 21.100 7.000 24.500 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END NAND2II

MACRO NAND2JJ
  CLASS CORE ;
  FOREIGN NAND2JJ 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
      RECT 16.400 11.500 17.400 14.900 ; # A|0.0@1
      RECT 6.000 13.900 17.400 14.900 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 14.900 ; # B|0.0@0
      RECT 11.200 6.700 12.200 12.500 ; # B|0.0@1
      RECT 21.600 6.700 22.600 12.500 ; # B|0.0@2
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 7.000 10.100 ; # Q|0.0@0
      RECT 16.400 9.100 20.000 10.100 ; # Q|0.0@1
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@2
      RECT 19.000 9.100 20.000 19.700 ; # Q|0.0@3
      RECT 3.400 18.700 20.000 19.700 ; # Q|0.0@4
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ;
      RECT 13.800 6.700 20.000 7.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 22.600 5.300 ;
      RECT 3.400 4.300 9.600 7.700 ;
      RECT 13.800 4.300 20.000 7.700 ;
      RECT 6.000 4.300 7.000 12.500 ;
      RECT 16.400 4.300 17.400 12.500 ;
      RECT 6.000 11.500 17.400 12.500 ;
      RECT 21.600 11.500 22.600 14.900 ;
      RECT 0.800 13.900 1.800 14.900 ;
      RECT 6.000 16.300 17.400 17.300 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 13.800 16.300 14.800 22.100 ;
      RECT 19.000 18.700 20.000 22.100 ;
      RECT 3.400 21.100 20.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 21.100 7.000 24.500 ;
      RECT 11.200 21.100 12.200 24.500 ;
      RECT 16.400 21.100 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END NAND2JJ

MACRO NAND3DD
  CLASS CORE ;
  FOREIGN NAND3DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 9.600 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 0.800 9.100 1.800 12.500 ;
      RECT 8.600 9.100 9.600 10.100 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END NAND3DD

MACRO NAND3EE
  CLASS CORE ;
  FOREIGN NAND3EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 9.600 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 9.100 9.600 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END NAND3EE

MACRO NAND3FF
  CLASS CORE ;
  FOREIGN NAND3FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # B|0.0@0
      RECT 6.000 13.900 9.600 14.900 ; # B|0.0@1
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 17.300 ; # C|0.0@0
      RECT 0.800 16.300 12.200 17.300 ; # C|0.0@1
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 14.800 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 14.800 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 7.700 ;
      RECT 8.600 9.100 12.200 12.500 ;
      RECT 3.400 11.500 12.200 12.500 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 11.200 9.100 12.200 14.900 ;
      RECT 3.400 18.700 12.200 22.100 ;
      RECT 3.400 21.100 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 6.000 4.300 14.800 5.300 ;
      RECT 6.000 4.300 7.000 7.700 ;
      RECT 8.600 9.100 12.200 12.500 ;
      RECT 0.800 11.500 12.200 12.500 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 11.200 9.100 12.200 14.900 ;
      RECT 3.400 18.700 12.200 22.100 ;
      RECT 3.400 21.100 14.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 18.700 7.000 24.500 ;
      RECT 11.200 18.700 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 14.800 29.300 ;
  END
END NAND3FF

MACRO NAND3GG
  CLASS CORE ;
  FOREIGN NAND3GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
      RECT 6.000 13.900 12.200 14.900 ; # B|0.0@1
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 22.100 ; # C|0.0@0
      RECT 16.400 13.900 17.400 22.100 ; # C|0.0@1
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 11.200 9.100 14.800 10.100 ; # Q|0.0@1
      RECT 13.800 9.100 14.800 17.300 ; # Q|0.0@2
      RECT 3.400 16.300 4.400 17.300 ; # Q|0.0@3
      RECT 8.600 16.300 9.600 17.300 ; # Q|0.0@4
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@5
      RECT 11.200 18.700 12.200 19.700 ; # Q|0.0@6
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 11.200 6.700 14.800 7.700 ;
      RECT 8.600 9.100 9.600 10.100 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 11.200 11.500 12.200 12.500 ;
      RECT 3.400 13.900 4.400 14.900 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 18.700 9.600 22.100 ;
      RECT 13.800 18.700 14.800 22.100 ;
      RECT 3.400 21.100 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 4.300 9.600 12.500 ;
      RECT 16.400 4.300 17.400 5.300 ;
      RECT 8.600 6.700 14.800 7.700 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 12.200 12.500 ;
      RECT 3.400 13.900 7.000 14.900 ;
      RECT 11.200 11.500 12.200 14.900 ;
      RECT 16.400 13.900 17.400 14.900 ;
      RECT 3.400 13.900 4.400 24.500 ;
      RECT 8.600 16.300 9.600 24.500 ;
      RECT 13.800 16.300 14.800 24.500 ;
      RECT 3.400 21.100 14.800 24.500 ;
      RECT 0.800 23.500 17.400 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NAND3GG

MACRO NAND3HH
  CLASS CORE ;
  FOREIGN NAND3HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 12.500 ; # A|0.0@0
      RECT 16.400 6.700 22.600 7.700 ; # A|0.0@1
      RECT 21.600 6.700 22.600 14.900 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 19.700 ; # Q|0.0@0
      RECT 8.600 9.100 14.800 10.100 ; # Q|0.0@1
      RECT 13.800 9.100 14.800 17.300 ; # Q|0.0@2
      RECT 3.400 18.700 7.000 19.700 ; # Q|0.0@3
      RECT 11.200 18.700 12.200 19.700 ; # Q|0.0@4
      RECT 16.400 18.700 17.400 19.700 ; # Q|0.0@5
      RECT 21.600 18.700 25.200 19.700 ; # Q|0.0@6
      RECT 3.400 18.700 4.400 22.100 ; # Q|0.0@7
      RECT 8.600 21.100 9.600 22.100 ; # Q|0.0@8
      RECT 13.800 21.100 14.800 22.100 ; # Q|0.0@9
      RECT 19.000 21.100 20.000 22.100 ; # Q|0.0@10
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 14.800 7.700 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 3.400 16.300 12.200 17.300 ;
      RECT 16.400 16.300 22.600 17.300 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 13.800 18.700 14.800 19.700 ;
      RECT 19.000 16.300 20.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 16.400 4.300 17.400 5.300 ;
      RECT 24.200 4.300 25.200 10.100 ;
      RECT 8.600 6.700 14.800 7.700 ;
      RECT 0.800 9.100 1.800 12.500 ;
      RECT 8.600 6.700 9.600 10.100 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 11.200 13.900 12.200 17.300 ;
      RECT 3.400 16.300 12.200 17.300 ;
      RECT 16.400 16.300 22.600 17.300 ;
      RECT 3.400 16.300 4.400 22.100 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 13.800 18.700 14.800 22.100 ;
      RECT 19.000 16.300 20.000 22.100 ;
      RECT 24.200 18.700 25.200 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END NAND3HH

MACRO NAND4CC
  CLASS CORE ;
  FOREIGN NAND4CC 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 12.200 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 21.100 4.400 22.100 ;
      RECT 8.600 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 8.600 9.100 12.200 10.100 ;
      RECT 8.600 9.100 9.600 12.500 ;
      RECT 0.800 13.900 7.000 14.900 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 18.700 9.600 22.100 ;
      RECT 8.600 21.100 12.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 21.100 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NAND4CC

MACRO NAND4DD
  CLASS CORE ;
  FOREIGN NAND4DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 12.200 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 21.100 4.400 22.100 ;
      RECT 8.600 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 11.200 9.100 12.200 10.100 ;
      RECT 8.600 11.500 9.600 12.500 ;
      RECT 0.800 13.900 7.000 14.900 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 18.700 9.600 22.100 ;
      RECT 8.600 21.100 12.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 21.100 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NAND4DD

MACRO NAND4FF
  CLASS CORE ;
  FOREIGN NAND4FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 20.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 21.600 4.300 22.600 5.300 ;
      RECT 11.200 9.100 12.200 10.100 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 8.600 13.900 9.600 22.100 ;
      RECT 13.800 13.900 14.800 22.100 ;
      RECT 3.400 13.900 4.400 22.100 ;
      RECT 19.000 16.300 20.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END NAND4FF

MACRO NAND4GG
  CLASS CORE ;
  FOREIGN NAND4GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 9.600 12.500 ; # B|0.0@0
      RECT 6.000 11.500 7.000 14.900 ; # B|0.0@1
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 12.500 ; # C|0.0@0
      RECT 19.000 6.700 20.000 12.500 ; # C|0.0@1
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 22.100 ; # D|0.0@0
      RECT 21.600 13.900 22.600 22.100 ; # D|0.0@1
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 17.400 10.100 ; # Q|0.0@0
      RECT 16.400 9.100 17.400 19.700 ; # Q|0.0@1
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@2
      RECT 11.200 18.700 12.200 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 17.400 7.700 ;
      RECT 8.600 6.700 12.200 10.100 ;
      RECT 11.200 11.500 14.800 12.500 ;
      RECT 3.400 13.900 4.400 22.100 ;
      RECT 13.800 11.500 14.800 22.100 ;
      RECT 19.000 13.900 20.000 22.100 ;
      RECT 8.600 16.300 14.800 17.300 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 3.400 21.100 20.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 19.000 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 22.600 5.300 ;
      RECT 6.000 4.300 17.400 7.700 ;
      RECT 8.600 4.300 12.200 12.500 ;
      RECT 6.000 11.500 14.800 12.500 ;
      RECT 19.000 11.500 22.600 17.300 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 13.800 11.500 14.800 24.500 ;
      RECT 3.400 13.900 4.400 24.500 ;
      RECT 8.600 16.300 14.800 17.300 ;
      RECT 8.600 16.300 9.600 24.500 ;
      RECT 19.000 11.500 20.000 24.500 ;
      RECT 3.400 21.100 20.000 24.500 ;
      RECT 0.800 23.500 22.600 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END NAND4GG

MACRO NAND4HH
  CLASS CORE ;
  FOREIGN NAND4HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 33.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 9.100 30.400 10.100 ; # B|0.0@0
      RECT 11.200 11.500 12.200 12.500 ; # B|0.0@1
      RECT 29.400 9.100 30.400 12.500 ; # B|0.0@2
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 11.500 25.200 12.500 ; # C|0.0@0
      RECT 6.000 13.900 7.000 14.900 ; # C|0.0@1
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 22.100 ; # D|0.0@0
      RECT 21.600 16.300 22.600 22.100 ; # D|0.0@1
      RECT 32.000 18.700 33.000 22.100 ; # D|0.0@2
      RECT 6.000 21.100 7.000 22.100 ; # D|0.0@3
      RECT 11.200 21.100 12.200 22.100 ; # D|0.0@4
      RECT 16.400 21.100 17.400 22.100 ; # D|0.0@5
      RECT 26.800 21.100 27.800 22.100 ; # D|0.0@6
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 33.000 7.700 ; # Q|0.0@1
      RECT 3.400 6.700 4.400 17.300 ; # Q|0.0@2
      RECT 11.200 9.100 12.200 10.100 ; # Q|0.0@3
      RECT 32.000 6.700 33.000 17.300 ; # Q|0.0@4
      RECT 29.400 16.300 33.000 17.300 ; # Q|0.0@5
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@6
      RECT 11.200 18.700 12.200 19.700 ; # Q|0.0@7
      RECT 16.400 18.700 17.400 19.700 ; # Q|0.0@8
      RECT 24.200 18.700 27.800 19.700 ; # Q|0.0@9
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 33.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 33.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 11.200 6.700 12.200 7.700 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 13.800 9.100 14.800 22.100 ;
      RECT 13.800 11.500 17.400 17.300 ;
      RECT 26.800 11.500 27.800 14.900 ;
      RECT 11.200 13.900 30.400 14.900 ;
      RECT 6.000 16.300 20.000 17.300 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 19.000 13.900 20.000 22.100 ;
      RECT 29.400 18.700 30.400 22.100 ;
      RECT 24.200 21.100 25.200 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 33.000 5.300 ;
      RECT 11.200 4.300 12.200 10.100 ;
      RECT 32.000 4.300 33.000 10.100 ;
      RECT 0.800 9.100 1.800 12.500 ;
      RECT 8.600 9.100 14.800 10.100 ;
      RECT 8.600 9.100 9.600 12.500 ;
      RECT 13.800 11.500 17.400 17.300 ;
      RECT 26.800 11.500 27.800 14.900 ;
      RECT 11.200 13.900 30.400 14.900 ;
      RECT 6.000 16.300 20.000 17.300 ;
      RECT 24.200 13.900 25.200 22.100 ;
      RECT 29.400 16.300 33.000 19.700 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 8.600 16.300 9.600 22.100 ;
      RECT 13.800 9.100 14.800 22.100 ;
      RECT 19.000 13.900 20.000 22.100 ;
      RECT 29.400 13.900 30.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 32.000 23.500 33.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
  END
END NAND4HH

MACRO NAND5FF
  CLASS CORE ;
  FOREIGN NAND5FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 12.500 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 9.100 25.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 20.000 7.700 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 16.400 6.700 20.000 19.700 ;
      RECT 16.400 11.500 22.600 19.700 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 13.900 22.600 14.900 ;
      RECT 8.600 13.900 12.200 19.700 ;
      RECT 3.400 18.700 22.600 19.700 ;
    LAYER cont2 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 8.600 4.300 12.200 7.700 ;
      RECT 6.000 6.700 25.200 7.700 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 16.400 6.700 25.200 10.100 ;
      RECT 16.400 6.700 22.600 19.700 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 8.600 13.900 22.600 19.700 ;
      RECT 3.400 16.300 25.200 19.700 ;
      RECT 3.400 13.900 4.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END NAND5FF

MACRO NAND6FF
  CLASS CORE ;
  FOREIGN NAND6FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # E|0.0@0
    END
  END E
  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 9.100 17.400 12.500 ; # F|0.0@0
    END
  END F
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 9.100 27.800 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 16.400 6.700 20.000 7.700 ;
      RECT 19.000 9.100 25.200 10.100 ;
      RECT 19.000 6.700 20.000 19.700 ;
      RECT 24.200 9.100 25.200 19.700 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 13.800 16.300 25.200 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 13.800 18.700 27.800 19.700 ;
    LAYER cont2 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 16.400 4.300 20.000 10.100 ;
      RECT 24.200 4.300 25.200 5.300 ;
      RECT 6.000 6.700 12.200 7.700 ;
      RECT 16.400 6.700 22.600 10.100 ;
      RECT 26.800 6.700 27.800 10.100 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 16.400 9.100 27.800 10.100 ;
      RECT 19.000 9.100 25.200 19.700 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 8.600 13.900 14.800 14.900 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 13.800 16.300 27.800 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 24.200 23.500 25.200 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END NAND6FF

MACRO NINVJJ
  CLASS CORE ;
  FOREIGN NINVJJ 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 19.700 ; # Q|0.0@0
      RECT 8.600 13.900 14.800 14.900 ; # Q|0.0@1
      RECT 8.600 13.900 9.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 10.700 21.600 12.300 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 16.400 6.700 17.400 10.100 ;
      RECT 3.400 6.700 9.600 12.500 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 0.800 16.300 7.000 19.700 ;
      RECT 0.800 16.300 4.400 22.100 ;
      RECT 11.200 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 11.200 4.300 12.200 12.500 ;
      RECT 0.800 6.700 17.400 7.700 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 16.400 6.700 17.400 10.100 ;
      RECT 3.400 6.700 12.200 12.500 ;
      RECT 3.400 6.700 7.000 19.700 ;
      RECT 0.800 16.300 14.800 17.300 ;
      RECT 0.800 16.300 9.600 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 0.800 16.300 4.400 22.100 ;
      RECT 8.600 21.100 12.200 24.500 ;
      RECT 0.800 16.300 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END NINVJJ

MACRO NINVKK
  CLASS CORE ;
  FOREIGN NINVKK 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 6.700 14.800 7.700 ; # Q|0.0@0
      RECT 21.600 6.700 25.200 7.700 ; # Q|0.0@1
      RECT 24.200 6.700 25.200 14.900 ; # Q|0.0@2
      RECT 11.200 13.900 25.200 14.900 ; # Q|0.0@3
      RECT 11.200 13.900 12.200 17.300 ; # Q|0.0@4
      RECT 16.400 13.900 17.400 19.700 ; # Q|0.0@5
      RECT 21.600 13.900 22.600 19.700 ; # Q|0.0@6
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.500 21.600 15.100 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 11.200 6.700 12.200 12.500 ;
      RECT 16.400 6.700 20.000 10.100 ;
      RECT 3.400 9.100 12.200 10.100 ;
      RECT 3.400 6.700 4.400 17.300 ;
      RECT 8.600 9.100 12.200 12.500 ;
      RECT 0.800 13.900 9.600 17.300 ;
      RECT 0.800 13.900 1.800 19.700 ;
      RECT 6.000 13.900 7.000 19.700 ;
      RECT 11.200 18.700 12.200 19.700 ;
      RECT 13.800 21.100 14.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 25.200 5.300 ;
      RECT 3.400 4.300 12.200 12.500 ;
      RECT 16.400 4.300 20.000 12.500 ;
      RECT 24.200 4.300 25.200 10.100 ;
      RECT 3.400 9.100 20.000 12.500 ;
      RECT 3.400 11.500 22.600 12.500 ;
      RECT 0.800 13.900 9.600 17.300 ;
      RECT 0.800 16.300 25.200 17.300 ;
      RECT 0.800 13.900 1.800 19.700 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 11.200 16.300 12.200 19.700 ;
      RECT 16.400 16.300 17.400 19.700 ;
      RECT 21.600 16.300 25.200 19.700 ;
      RECT 13.800 21.100 14.800 24.500 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END NINVKK

MACRO NOR2DD
  CLASS CORE ;
  FOREIGN NOR2DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@0
      RECT 3.400 18.700 7.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 16.300 7.000 17.300 ;
    LAYER cont2 ;
      RECT 0.800 4.300 7.000 5.300 ;
      RECT 3.400 9.100 4.400 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 7.000 12.500 ;
      RECT 6.000 16.300 7.000 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END NOR2DD

MACRO NOR2FF
  CLASS CORE ;
  FOREIGN NOR2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 14.900 ; # B|0.0@0
      RECT 8.600 6.700 12.200 7.700 ; # B|0.0@1
      RECT 11.200 6.700 12.200 12.500 ; # B|0.0@2
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 7.000 10.100 ;
      RECT 8.600 11.500 9.600 12.500 ;
    LAYER cont2 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 8.600 4.300 9.600 5.300 ;
      RECT 6.000 6.700 7.000 10.100 ;
      RECT 6.000 9.100 9.600 10.100 ;
      RECT 3.400 11.500 4.400 12.500 ;
      RECT 8.600 11.500 12.200 12.500 ;
      RECT 11.200 11.500 12.200 14.900 ;
      RECT 6.000 16.300 7.000 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NOR2FF

MACRO NOR2GG
  CLASS CORE ;
  FOREIGN NOR2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 7.000 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # B|0.0@0
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@1
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 14.800 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 14.800 17.300 ; # Q|0.0@1
      RECT 8.600 16.300 14.800 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 3.400 11.500 7.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 3.400 4.300 7.000 7.700 ;
      RECT 11.200 4.300 12.200 7.700 ;
      RECT 6.000 9.100 9.600 14.900 ;
      RECT 0.800 11.500 9.600 12.500 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 3.400 11.500 7.000 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 3.400 18.700 14.800 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NOR2GG

MACRO NOR2HH
  CLASS CORE ;
  FOREIGN NOR2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 14.800 10.100 ; # A|0.0@0
      RECT 6.000 11.500 7.000 12.500 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 19.700 ; # B|0.0@0
      RECT 11.200 11.500 12.200 19.700 ; # B|0.0@1
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 16.400 6.700 17.400 17.300 ; # Q|0.0@1
      RECT 3.400 9.100 4.400 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 11.200 6.700 14.800 7.700 ;
      RECT 6.000 6.700 7.000 10.100 ;
      RECT 6.000 13.900 7.000 22.100 ;
      RECT 3.400 18.700 9.600 22.100 ;
      RECT 16.400 18.700 17.400 19.700 ;
      RECT 0.800 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 17.400 5.300 ;
      RECT 0.800 4.300 7.000 7.700 ;
      RECT 11.200 4.300 14.800 7.700 ;
      RECT 6.000 4.300 7.000 10.100 ;
      RECT 13.800 4.300 14.800 14.900 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 13.900 7.000 22.100 ;
      RECT 11.200 13.900 14.800 14.900 ;
      RECT 16.400 16.300 17.400 19.700 ;
      RECT 3.400 18.700 9.600 22.100 ;
      RECT 0.800 21.100 12.200 22.100 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 11.200 21.100 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END NOR2HH

MACRO NOR3DD
  CLASS CORE ;
  FOREIGN NOR3DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 14.800 10.100 ; # Q|0.0@0
      RECT 6.000 9.100 7.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 4.300 4.400 5.300 ;
      RECT 11.200 4.300 12.200 7.700 ;
      RECT 6.000 6.700 14.800 7.700 ;
      RECT 3.400 9.100 7.000 10.100 ;
      RECT 13.800 6.700 14.800 12.500 ;
      RECT 3.400 9.100 4.400 12.500 ;
      RECT 8.600 11.500 14.800 12.500 ;
      RECT 0.800 13.900 1.800 14.900 ;
      RECT 8.600 11.500 9.600 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
  END
END NOR3DD

MACRO NOR3FF
  CLASS CORE ;
  FOREIGN NOR3FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 17.400 10.100 ; # A|0.0@0
      RECT 19.000 11.500 20.000 12.500 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # C|0.0@0
      RECT 0.800 13.900 4.400 14.900 ; # C|0.0@1
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 12.200 7.700 ; # Q|0.0@0
      RECT 16.400 6.700 17.400 7.700 ; # Q|0.0@1
      RECT 21.600 6.700 22.600 19.700 ; # Q|0.0@2
      RECT 8.600 18.700 22.600 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 12.500 ;
      RECT 13.800 6.700 14.800 7.700 ;
      RECT 19.000 6.700 20.000 10.100 ;
      RECT 3.400 9.100 12.200 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 9.100 12.200 17.300 ;
      RECT 6.000 13.900 12.200 17.300 ;
      RECT 6.000 16.300 20.000 17.300 ;
      RECT 6.000 6.700 7.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 22.600 5.300 ;
      RECT 3.400 4.300 7.000 14.900 ;
      RECT 13.800 4.300 14.800 7.700 ;
      RECT 19.000 4.300 20.000 10.100 ;
      RECT 3.400 9.100 12.200 10.100 ;
      RECT 0.800 11.500 7.000 14.900 ;
      RECT 11.200 9.100 12.200 17.300 ;
      RECT 0.800 13.900 14.800 14.900 ;
      RECT 6.000 16.300 22.600 17.300 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 21.600 16.300 22.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
  END
END NOR3FF

MACRO NOR3GG
  CLASS CORE ;
  FOREIGN NOR3GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # A|0.0@0
      RECT 21.600 11.500 22.600 12.500 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 7.000 10.100 ; # B|0.0@0
      RECT 19.000 9.100 20.000 10.100 ; # B|0.0@1
      RECT 3.400 9.100 4.400 12.500 ; # B|0.0@2
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 11.500 27.800 22.100 ; # C|0.0@0
      RECT 0.800 13.900 1.800 22.100 ; # C|0.0@1
      RECT 0.800 21.100 4.400 22.100 ; # C|0.0@2
      RECT 11.200 21.100 17.400 22.100 ; # C|0.0@3
      RECT 24.200 21.100 27.800 22.100 ; # C|0.0@4
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 13.800 6.700 17.400 7.700 ; # Q|0.0@1
      RECT 21.600 6.700 25.200 7.700 ; # Q|0.0@2
      RECT 24.200 6.700 25.200 17.300 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 7.700 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 19.000 6.700 20.000 7.700 ;
      RECT 8.600 9.100 17.400 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 11.200 11.500 20.000 19.700 ;
      RECT 8.600 13.900 22.600 19.700 ;
      RECT 6.000 16.300 22.600 19.700 ;
      RECT 6.000 18.700 25.200 19.700 ;
      RECT 6.000 16.300 9.600 22.100 ;
      RECT 19.000 13.900 22.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 17.400 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 25.200 5.300 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 11.200 4.300 12.200 19.700 ;
      RECT 19.000 4.300 20.000 22.100 ;
      RECT 8.600 9.100 20.000 19.700 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 8.600 13.900 22.600 19.700 ;
      RECT 26.800 13.900 27.800 14.900 ;
      RECT 6.000 16.300 22.600 19.700 ;
      RECT 6.000 18.700 25.200 19.700 ;
      RECT 6.000 16.300 9.600 22.100 ;
      RECT 19.000 13.900 22.600 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END NOR3GG

MACRO NOR3HH
  CLASS CORE ;
  FOREIGN NOR3HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 44.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 9.100 35.600 10.100 ; # A|0.0@0
      RECT 19.000 11.500 20.000 12.500 ; # A|0.0@1
      RECT 34.600 9.100 35.600 14.900 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 11.500 30.400 22.100 ; # C|0.0@0
      RECT 0.800 13.900 1.800 22.100 ; # C|0.0@1
      RECT 42.400 13.900 43.400 22.100 ; # C|0.0@2
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 12.200 7.700 ; # Q|0.0@0
      RECT 16.400 6.700 17.400 7.700 ; # Q|0.0@1
      RECT 37.200 6.700 43.400 7.700 ; # Q|0.0@2
      RECT 6.000 9.100 7.000 19.700 ; # Q|0.0@3
      RECT 39.800 6.700 40.800 17.300 ; # Q|0.0@4
      RECT 6.000 16.300 9.600 19.700 ; # Q|0.0@5
      RECT 34.600 16.300 40.800 17.300 ; # Q|0.0@6
      RECT 34.600 16.300 35.600 19.700 ; # Q|0.0@7
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 44.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 44.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 13.800 6.700 14.800 22.100 ;
      RECT 19.000 6.700 35.600 7.700 ;
      RECT 8.600 9.100 27.800 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 8.600 9.100 17.400 14.900 ;
      RECT 21.600 6.700 27.800 22.100 ;
      RECT 42.400 11.500 43.400 12.500 ;
      RECT 8.600 13.900 27.800 14.900 ;
      RECT 13.800 13.900 27.800 22.100 ;
      RECT 3.400 21.100 27.800 22.100 ;
      RECT 32.000 21.100 40.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 39.800 -0.500 40.800 0.500 ;
      RECT 0.800 4.300 43.400 5.300 ;
      RECT 3.400 4.300 7.000 7.700 ;
      RECT 13.800 4.300 14.800 24.500 ;
      RECT 19.000 4.300 35.600 7.700 ;
      RECT 42.400 4.300 43.400 7.700 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 8.600 9.100 27.800 10.100 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 8.600 9.100 17.400 14.900 ;
      RECT 21.600 4.300 27.800 24.500 ;
      RECT 42.400 11.500 43.400 14.900 ;
      RECT 8.600 13.900 30.400 14.900 ;
      RECT 34.600 13.900 38.200 14.900 ;
      RECT 8.600 9.100 9.600 24.500 ;
      RECT 13.800 13.900 27.800 24.500 ;
      RECT 34.600 13.900 35.600 24.500 ;
      RECT 34.600 18.700 40.800 24.500 ;
      RECT 3.400 21.100 27.800 24.500 ;
      RECT 32.000 21.100 40.800 24.500 ;
      RECT 0.800 23.500 43.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
  END
END NOR3HH

MACRO NOR4DD
  CLASS CORE ;
  FOREIGN NOR4DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 20.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 19.700 ; # B|0.0@0
      RECT 13.800 11.500 14.800 19.700 ; # B|0.0@1
      RECT 6.000 18.700 14.800 19.700 ; # B|0.0@2
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 9.100 17.400 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 6.700 9.600 7.700 ; # Q|0.0@0
      RECT 11.200 9.100 12.200 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 18.100 16.800 19.800 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 20.800 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 20.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 7.700 ;
      RECT 11.200 6.700 14.800 7.700 ;
      RECT 13.800 6.700 14.800 10.100 ;
      RECT 8.600 11.500 9.600 17.300 ;
      RECT 16.400 13.900 17.400 22.100 ;
      RECT 16.400 16.300 20.000 17.300 ;
    LAYER cont2 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 3.400 4.300 7.000 7.700 ;
      RECT 11.200 4.300 14.800 7.700 ;
      RECT 13.800 4.300 14.800 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 9.600 12.500 ;
      RECT 16.400 11.500 17.400 24.500 ;
      RECT 8.600 11.500 9.600 17.300 ;
      RECT 16.400 16.300 20.000 24.500 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END NOR4DD

MACRO NOR4FF
  CLASS CORE ;
  FOREIGN NOR4FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 33.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 17.300 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 7.700 ; # Q|0.0@0
      RECT 0.800 11.500 1.800 19.700 ; # Q|0.0@1
      RECT 0.800 18.700 20.000 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 33.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 33.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 16.400 6.700 22.600 17.300 ;
      RECT 0.800 9.100 22.600 10.100 ;
      RECT 3.400 6.700 4.400 12.500 ;
      RECT 8.600 9.100 22.600 12.500 ;
      RECT 11.200 6.700 12.200 17.300 ;
      RECT 6.000 16.300 22.600 17.300 ;
      RECT 21.600 6.700 22.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 14.800 10.100 ;
      RECT 0.800 6.700 22.600 10.100 ;
      RECT 0.800 4.300 4.400 12.500 ;
      RECT 8.600 6.700 22.600 12.500 ;
      RECT 11.200 4.300 12.200 22.100 ;
      RECT 16.400 6.700 22.600 22.100 ;
      RECT 6.000 16.300 22.600 17.300 ;
      RECT 0.800 21.100 22.600 22.100 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 19.000 6.700 20.000 24.500 ;
      RECT 32.000 23.500 33.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
  END
END NOR4FF

MACRO NOR4GG
  CLASS CORE ;
  FOREIGN NOR4GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 41.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 9.100 27.800 14.900 ; # A|0.0@0
      RECT 11.200 13.900 12.200 14.900 ; # A|0.0@1
      RECT 16.400 13.900 27.800 14.900 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 6.700 20.000 12.500 ; # B|0.0@0
      RECT 32.000 6.700 33.000 7.700 ; # B|0.0@1
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@2
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 7.700 ; # C|0.0@0
      RECT 11.200 9.100 14.800 10.100 ; # C|0.0@1
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 17.300 ; # D|0.0@0
      RECT 3.400 16.300 9.600 17.300 ; # D|0.0@1
      RECT 13.800 16.300 14.800 17.300 ; # D|0.0@2
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
      RECT 6.000 6.700 9.600 7.700 ; # Q|0.0@1
      RECT 0.800 18.700 9.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 37.100 15.600 39.000 23.600 ; # VDD|0.0@0
      RECT 0.000 23.600 41.600 29.200 ; # VDD|0.0@1
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 41.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 11.200 6.700 12.200 7.700 ;
      RECT 21.600 6.700 30.400 7.700 ;
      RECT 3.400 9.100 9.600 10.100 ;
      RECT 16.400 9.100 17.400 12.500 ;
      RECT 29.400 6.700 30.400 10.100 ;
      RECT 6.000 9.100 7.000 12.500 ;
      RECT 11.200 11.500 17.400 12.500 ;
      RECT 13.800 11.500 14.800 14.900 ;
      RECT 37.200 13.900 40.800 14.900 ;
      RECT 11.200 16.300 12.200 22.100 ;
      RECT 16.400 16.300 20.000 22.100 ;
      RECT 39.800 13.900 40.800 22.100 ;
      RECT 11.200 18.700 30.400 22.100 ;
      RECT 0.800 21.100 30.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 37.200 -0.500 40.800 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 19.000 4.300 33.000 5.300 ;
      RECT 37.200 4.300 40.800 5.300 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 11.200 4.300 12.200 7.700 ;
      RECT 21.600 4.300 33.000 7.700 ;
      RECT 3.400 9.100 9.600 10.100 ;
      RECT 13.800 9.100 17.400 12.500 ;
      RECT 29.400 4.300 30.400 10.100 ;
      RECT 6.000 11.500 17.400 12.500 ;
      RECT 8.600 11.500 14.800 14.900 ;
      RECT 37.200 13.900 40.800 17.300 ;
      RECT 11.200 11.500 12.200 22.100 ;
      RECT 16.400 16.300 20.000 22.100 ;
      RECT 11.200 18.700 30.400 22.100 ;
      RECT 39.800 13.900 40.800 24.500 ;
      RECT 0.800 21.100 30.400 22.100 ;
      RECT 37.200 21.100 40.800 24.500 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 26.800 18.700 30.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
  END
END NOR4GG

MACRO NOR4HH
  CLASS CORE ;
  FOREIGN NOR4HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 59.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 11.500 33.000 14.900 ; # A|0.0@0
      RECT 11.200 13.900 14.800 14.900 ; # A|0.0@1
      RECT 21.600 13.900 27.800 14.900 ; # A|0.0@2
      RECT 32.000 13.900 38.200 14.900 ; # A|0.0@3
      RECT 45.000 13.900 48.600 14.900 ; # A|0.0@4
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 34.600 9.100 35.600 12.500 ; # B|0.0@0
      RECT 8.600 11.500 9.600 12.500 ; # B|0.0@1
      RECT 19.000 11.500 20.000 12.500 ; # B|0.0@2
      RECT 50.200 11.500 51.200 12.500 ; # B|0.0@3
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 39.800 6.700 43.400 7.700 ; # C|0.0@0
      RECT 11.200 9.100 12.200 10.100 ; # C|0.0@1
      RECT 16.400 9.100 17.400 10.100 ; # C|0.0@2
      RECT 52.800 11.500 53.800 12.500 ; # C|0.0@3
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # D|0.0@0
      RECT 55.400 11.500 56.400 14.900 ; # D|0.0@1
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
      RECT 58.000 6.700 59.000 19.700 ; # Q|0.0@1
      RECT 0.800 18.700 59.000 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 59.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 59.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 21.600 6.700 38.200 7.700 ;
      RECT 47.600 6.700 56.400 10.100 ;
      RECT 3.400 6.700 9.600 10.100 ;
      RECT 13.800 9.100 14.800 12.500 ;
      RECT 21.600 6.700 25.200 12.500 ;
      RECT 29.400 6.700 33.000 10.100 ;
      RECT 42.400 9.100 56.400 10.100 ;
      RECT 6.000 6.700 7.000 12.500 ;
      RECT 11.200 11.500 17.400 12.500 ;
      RECT 29.400 6.700 30.400 17.300 ;
      RECT 37.200 11.500 48.600 12.500 ;
      RECT 16.400 13.900 20.000 17.300 ;
      RECT 39.800 11.500 43.400 17.300 ;
      RECT 3.400 16.300 56.400 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 13.800 -0.500 17.400 0.500 ;
      RECT 39.800 -0.500 46.000 0.500 ;
      RECT 52.800 -0.500 53.800 0.500 ;
      RECT 58.000 -0.500 59.000 0.500 ;
      RECT 0.800 4.300 17.400 5.300 ;
      RECT 21.600 4.300 59.000 5.300 ;
      RECT 3.400 4.300 17.400 7.700 ;
      RECT 21.600 4.300 38.200 7.700 ;
      RECT 45.000 4.300 56.400 10.100 ;
      RECT 3.400 4.300 9.600 10.100 ;
      RECT 13.800 4.300 17.400 12.500 ;
      RECT 21.600 4.300 25.200 12.500 ;
      RECT 29.400 4.300 33.000 10.100 ;
      RECT 37.200 9.100 56.400 10.100 ;
      RECT 6.000 11.500 30.400 12.500 ;
      RECT 37.200 9.100 51.200 12.500 ;
      RECT 8.600 11.500 12.200 17.300 ;
      RECT 16.400 11.500 20.000 17.300 ;
      RECT 29.400 4.300 30.400 19.700 ;
      RECT 39.800 9.100 43.400 17.300 ;
      RECT 47.600 4.300 51.200 17.300 ;
      RECT 3.400 16.300 56.400 17.300 ;
      RECT 11.200 11.500 12.200 19.700 ;
      RECT 47.600 4.300 48.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 19.000 23.500 22.600 24.500 ;
      RECT 39.800 23.500 40.800 24.500 ;
      RECT 58.000 23.500 59.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 19.000 28.300 22.600 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
  END
END NOR4HH

MACRO NOR5FF
  CLASS CORE ;
  FOREIGN NOR5FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 26.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 25.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 26.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 26.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 20.000 7.700 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 16.400 9.100 22.600 19.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 13.800 16.300 22.600 19.700 ;
      RECT 6.000 18.700 22.600 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 19.000 4.300 25.200 7.700 ;
      RECT 3.400 6.700 25.200 7.700 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 16.400 6.700 22.600 19.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 0.800 13.900 1.800 14.900 ;
      RECT 13.800 13.900 22.600 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 13.800 16.300 25.200 19.700 ;
      RECT 6.000 18.700 25.200 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 19.000 28.300 22.600 29.300 ;
  END
END NOR5FF

MACRO NOR6FF
  CLASS CORE ;
  FOREIGN NOR6FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 11.500 17.400 14.900 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 12.500 ; # E|0.0@0
    END
  END E
  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # F|0.0@0
    END
  END F
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 6.700 27.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 25.200 7.700 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 19.000 6.700 25.200 22.100 ;
      RECT 8.600 6.700 12.200 12.500 ;
      RECT 8.600 6.700 9.600 22.100 ;
      RECT 16.400 16.300 25.200 22.100 ;
      RECT 8.600 18.700 25.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 16.400 4.300 17.400 7.700 ;
      RECT 21.600 4.300 27.800 7.700 ;
      RECT 3.400 6.700 27.800 7.700 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 19.000 6.700 25.200 22.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 8.600 11.500 14.800 12.500 ;
      RECT 8.600 6.700 9.600 22.100 ;
      RECT 13.800 13.900 25.200 14.900 ;
      RECT 16.400 16.300 27.800 19.700 ;
      RECT 8.600 18.700 27.800 19.700 ;
      RECT 8.600 18.700 25.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 18.700 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
  END
END NOR6FF

MACRO NTRIZKK
  CLASS CORE ;
  FOREIGN NTRIZKK 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 44.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 14.800 14.900 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 13.900 20.000 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 6.700 33.000 7.700 ; # Q|0.0@0
      RECT 37.200 6.700 38.200 7.700 ; # Q|0.0@1
      RECT 42.400 6.700 43.400 19.700 ; # Q|0.0@2
      RECT 29.400 18.700 30.400 19.700 ; # Q|0.0@3
      RECT 37.200 18.700 38.200 19.700 ; # Q|0.0@4
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 44.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 44.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ;
      RECT 11.200 6.700 30.400 7.700 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 39.800 6.700 40.800 22.100 ;
      RECT 8.600 9.100 9.600 12.500 ;
      RECT 13.800 9.100 40.800 10.100 ;
      RECT 0.800 11.500 9.600 12.500 ;
      RECT 21.600 9.100 40.800 17.300 ;
      RECT 6.000 16.300 40.800 17.300 ;
      RECT 6.000 16.300 27.800 19.700 ;
      RECT 32.000 9.100 35.600 22.100 ;
      RECT 8.600 21.100 40.800 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 26.800 -0.500 27.800 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 42.400 -0.500 43.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 11.200 4.300 43.400 5.300 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 11.200 4.300 17.400 10.100 ;
      RECT 21.600 4.300 22.600 19.700 ;
      RECT 26.800 4.300 30.400 17.300 ;
      RECT 34.600 4.300 35.600 22.100 ;
      RECT 39.800 4.300 40.800 10.100 ;
      RECT 0.800 9.100 17.400 10.100 ;
      RECT 21.600 9.100 40.800 10.100 ;
      RECT 3.400 9.100 14.800 12.500 ;
      RECT 21.600 9.100 38.200 17.300 ;
      RECT 3.400 9.100 4.400 17.300 ;
      RECT 13.800 4.300 14.800 17.300 ;
      RECT 21.600 13.900 40.800 17.300 ;
      RECT 3.400 16.300 40.800 17.300 ;
      RECT 0.800 18.700 1.800 19.700 ;
      RECT 6.000 16.300 7.000 19.700 ;
      RECT 11.200 16.300 12.200 19.700 ;
      RECT 16.400 16.300 17.400 19.700 ;
      RECT 21.600 9.100 27.800 19.700 ;
      RECT 32.000 9.100 35.600 22.100 ;
      RECT 39.800 13.900 40.800 22.100 ;
      RECT 8.600 21.100 9.600 24.500 ;
      RECT 26.800 21.100 43.400 22.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 8.600 23.500 25.200 24.500 ;
      RECT 29.400 21.100 30.400 24.500 ;
      RECT 37.200 21.100 38.200 24.500 ;
      RECT 42.400 21.100 43.400 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 29.400 28.300 30.400 29.300 ;
      RECT 37.200 28.300 38.200 29.300 ;
      RECT 42.400 28.300 43.400 29.300 ;
  END
END NTRIZKK

MACRO OAI211DD
  CLASS CORE ;
  FOREIGN OAI211DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 10.100 ; # Q|0.0@0
      RECT 0.800 9.100 4.400 10.100 ; # Q|0.0@1
      RECT 3.400 9.100 4.400 17.300 ; # Q|0.0@2
      RECT 6.000 18.700 12.200 19.700 ; # Q|0.0@3
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 6.000 6.700 9.600 10.100 ;
      RECT 8.600 6.700 9.600 12.500 ;
      RECT 6.000 13.900 7.000 17.300 ;
      RECT 11.200 16.300 12.200 17.300 ;
      RECT 3.400 18.700 4.400 19.700 ;
    LAYER cont2 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 3.400 4.300 12.200 7.700 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 0.800 6.700 1.800 12.500 ;
      RECT 6.000 4.300 9.600 12.500 ;
      RECT 6.000 11.500 14.800 12.500 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 3.400 16.300 7.000 19.700 ;
      RECT 11.200 16.300 14.800 19.700 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
  END
END OAI211DD

MACRO OAI211FF
  CLASS CORE ;
  FOREIGN OAI211FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # A|0.0@0
      RECT 11.200 11.500 12.200 12.500 ; # A|0.0@1
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 17.400 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 12.500 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
      RECT 21.600 16.300 22.600 19.700 ; # Q|0.0@1
      RECT 0.800 18.700 22.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 20.000 7.700 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 6.000 6.700 9.600 12.500 ;
      RECT 8.600 13.900 12.200 17.300 ;
      RECT 21.600 13.900 22.600 14.900 ;
      RECT 16.400 16.300 17.400 17.300 ;
    LAYER cont2 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 3.400 4.300 20.000 10.100 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 3.400 4.300 9.600 12.500 ;
      RECT 13.800 4.300 14.800 14.900 ;
      RECT 6.000 13.900 17.400 14.900 ;
      RECT 21.600 13.900 22.600 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 8.600 13.900 12.200 19.700 ;
      RECT 16.400 13.900 17.400 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END OAI211FF

MACRO OAI21DD
  CLASS CORE ;
  FOREIGN OAI21DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 12.500 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 4.400 7.700 ; # Q|0.0@0
      RECT 3.400 6.700 4.400 17.300 ; # Q|0.0@1
      RECT 3.400 16.300 7.000 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 9.600 7.700 ;
      RECT 8.600 16.300 9.600 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 9.600 5.300 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 9.600 7.700 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 6.000 11.500 9.600 19.700 ;
      RECT 3.400 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
  END
END OAI21DD

MACRO OAI21FF
  CLASS CORE ;
  FOREIGN OAI21FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # B|0.0@0
      RECT 8.600 13.900 9.600 14.900 ; # B|0.0@1
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 6.700 14.800 17.300 ; # Q|0.0@0
      RECT 6.000 16.300 7.000 17.300 ; # Q|0.0@1
      RECT 11.200 16.300 14.800 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 0.800 6.700 9.600 10.100 ;
      RECT 3.400 13.900 7.000 14.900 ;
      RECT 3.400 13.900 4.400 17.300 ;
      RECT 8.600 16.300 9.600 17.300 ;
    LAYER cont2 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 3.400 4.300 14.800 5.300 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 0.800 6.700 1.800 12.500 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 11.200 4.300 12.200 12.500 ;
      RECT 3.400 13.900 9.600 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 3.400 18.700 14.800 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END OAI21FF

MACRO OAI221DD
  CLASS CORE ;
  FOREIGN OAI221DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 16.300 9.600 17.300 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 16.300 7.000 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 13.900 1.800 17.300 ; # C|0.0@0
      RECT 11.200 16.300 12.200 17.300 ; # C|0.0@1
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 16.300 4.400 17.300 ; # D|0.0@0
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 16.300 17.400 17.300 ; # E|0.0@0
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 12.500 ; # Q|0.0@0
      RECT 13.800 16.300 14.800 22.100 ; # Q|0.0@1
      RECT 0.800 21.100 14.800 22.100 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 14.800 14.900 ;
      RECT 0.800 9.100 14.800 12.500 ;
      RECT 3.400 13.900 17.400 14.900 ;
      RECT 0.800 18.700 12.200 19.700 ;
    LAYER cont2 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 3.400 4.300 17.400 5.300 ;
      RECT 3.400 4.300 14.800 14.900 ;
      RECT 0.800 9.100 14.800 14.900 ;
      RECT 0.800 11.500 17.400 14.900 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 0.800 18.700 1.800 22.100 ;
      RECT 13.800 18.700 14.800 22.100 ;
      RECT 6.000 23.500 9.600 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OAI221DD

MACRO OAI22DD
  CLASS CORE ;
  FOREIGN OAI22DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 16.300 4.400 17.300 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 13.900 1.800 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 12.500 ; # C|0.0@0
      RECT 6.000 13.900 7.000 14.900 ; # C|0.0@1
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 17.300 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 9.600 10.100 ; # Q|0.0@0
      RECT 8.600 9.100 9.600 19.700 ; # Q|0.0@1
      RECT 6.000 18.700 9.600 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 10.100 ;
      RECT 3.400 11.500 7.000 12.500 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 6.000 16.300 7.000 17.300 ;
      RECT 11.200 18.700 12.200 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 8.600 6.700 12.200 10.100 ;
      RECT 3.400 11.500 7.000 12.500 ;
      RECT 11.200 6.700 12.200 12.500 ;
      RECT 0.800 13.900 4.400 14.900 ;
      RECT 6.000 16.300 7.000 19.700 ;
      RECT 11.200 16.300 12.200 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END OAI22DD

MACRO OAI22FF
  CLASS CORE ;
  FOREIGN OAI22FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 20.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 10.100 ; # A|0.0@0
      RECT 3.400 13.900 4.400 14.900 ; # A|0.0@1
      RECT 8.600 13.900 9.600 14.900 ; # A|0.0@2
      RECT 16.400 13.900 17.400 14.900 ; # A|0.0@3
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 20.000 10.100 ; # Q|0.0@0
      RECT 19.000 9.100 20.000 19.700 ; # Q|0.0@1
      RECT 6.000 18.700 20.000 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 20.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 20.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 14.800 7.700 ;
      RECT 8.600 6.700 12.200 10.100 ;
      RECT 3.400 11.500 4.400 12.500 ;
      RECT 8.600 6.700 9.600 12.500 ;
      RECT 16.400 11.500 17.400 12.500 ;
      RECT 3.400 16.300 17.400 17.300 ;
      RECT 3.400 16.300 4.400 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 3.400 4.300 17.400 5.300 ;
      RECT 6.000 6.700 20.000 7.700 ;
      RECT 8.600 4.300 12.200 12.500 ;
      RECT 0.800 11.500 12.200 12.500 ;
      RECT 16.400 11.500 17.400 17.300 ;
      RECT 3.400 16.300 17.400 17.300 ;
      RECT 3.400 16.300 7.000 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 23.500 12.200 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 12.200 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END OAI22FF

MACRO OAOIFF
  CLASS CORE ;
  FOREIGN OAOIFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 28.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 17.400 10.100 ; # A|0.0@0
      RECT 11.200 11.500 12.200 12.500 ; # A|0.0@1
      RECT 16.400 9.100 17.400 12.500 ; # A|0.0@2
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 9.600 10.100 ; # C|0.0@0
      RECT 0.800 9.100 1.800 12.500 ; # C|0.0@1
      RECT 8.600 9.100 9.600 12.500 ; # C|0.0@2
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 9.100 22.600 10.100 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 6.700 27.800 7.700 ; # Q|0.0@0
      RECT 26.800 6.700 27.800 19.700 ; # Q|0.0@1
      RECT 24.200 18.700 27.800 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 28.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 28.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 6.000 6.700 22.600 7.700 ;
      RECT 11.200 6.700 12.200 10.100 ;
      RECT 21.600 11.500 25.200 17.300 ;
      RECT 8.600 13.900 25.200 17.300 ;
      RECT 3.400 16.300 25.200 17.300 ;
      RECT 3.400 16.300 22.600 19.700 ;
      RECT 19.000 21.100 27.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 6.000 4.300 27.800 5.300 ;
      RECT 6.000 4.300 22.600 7.700 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 11.200 4.300 12.200 10.100 ;
      RECT 21.600 4.300 22.600 22.100 ;
      RECT 16.400 11.500 25.200 17.300 ;
      RECT 6.000 13.900 25.200 17.300 ;
      RECT 3.400 16.300 27.800 17.300 ;
      RECT 3.400 16.300 22.600 22.100 ;
      RECT 26.800 16.300 27.800 22.100 ;
      RECT 3.400 21.100 27.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 13.900 9.600 24.500 ;
      RECT 16.400 11.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OAOIFF

MACRO OR2EE
  CLASS CORE ;
  FOREIGN OR2EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 7.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 4.400 7.700 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 3.400 28.300 7.000 29.300 ;
  END
END OR2EE

MACRO OR2FF
  CLASS CORE ;
  FOREIGN OR2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 10.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 6.700 9.600 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 10.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 10.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 7.700 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 7.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 4.400 7.700 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 0.800 4.300 1.800 12.500 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 6.000 16.300 9.600 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 3.400 28.300 7.000 29.300 ;
  END
END OR2FF

MACRO OR2GG
  CLASS CORE ;
  FOREIGN OR2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 6.700 12.200 17.300 ; # Q|0.0@0
      RECT 8.600 18.700 9.600 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 7.000 7.700 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 6.000 11.500 9.600 17.300 ;
      RECT 0.800 13.900 1.800 19.700 ;
      RECT 0.800 16.300 9.600 17.300 ;
      RECT 0.800 16.300 7.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 12.200 5.300 ;
      RECT 0.800 4.300 7.000 7.700 ;
      RECT 11.200 4.300 12.200 10.100 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 3.400 11.500 9.600 12.500 ;
      RECT 0.800 13.900 1.800 19.700 ;
      RECT 6.000 11.500 9.600 19.700 ;
      RECT 0.800 16.300 9.600 19.700 ;
      RECT 0.800 18.700 12.200 19.700 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END OR2GG

MACRO OR2HH
  CLASS CORE ;
  FOREIGN OR2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 19.700 ; # B|0.0@0
      RECT 8.600 13.900 9.600 19.700 ; # B|0.0@1
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 9.100 17.400 17.300 ; # Q|0.0@0
      RECT 13.800 16.300 17.400 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 12.500 ;
      RECT 11.200 6.700 17.400 7.700 ;
      RECT 11.200 6.700 14.800 12.500 ;
      RECT 3.400 11.500 14.800 12.500 ;
      RECT 6.000 6.700 7.000 19.700 ;
      RECT 13.800 6.700 14.800 14.900 ;
      RECT 3.400 16.300 7.000 19.700 ;
      RECT 13.800 18.700 14.800 19.700 ;
    LAYER cont2 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 0.800 4.300 17.400 5.300 ;
      RECT 3.400 4.300 7.000 12.500 ;
      RECT 11.200 4.300 17.400 7.700 ;
      RECT 11.200 4.300 14.800 19.700 ;
      RECT 0.800 11.500 14.800 12.500 ;
      RECT 6.000 11.500 14.800 14.900 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 0.800 21.100 9.600 22.100 ;
      RECT 0.800 21.100 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
      RECT 8.600 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OR2HH

MACRO OR3EE
  CLASS CORE ;
  FOREIGN OR3EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 13.900 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 6.700 12.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 11.200 21.100 12.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 4.300 12.200 7.700 ;
      RECT 3.400 4.300 9.600 12.500 ;
      RECT 0.800 11.500 9.600 12.500 ;
      RECT 8.600 4.300 9.600 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 8.600 16.300 12.200 19.700 ;
      RECT 0.800 18.700 12.200 19.700 ;
      RECT 11.200 16.300 12.200 22.100 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 3.400 28.300 9.600 29.300 ;
  END
END OR3EE

MACRO OR3FF
  CLASS CORE ;
  FOREIGN OR3FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 9.100 12.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
    LAYER cont2 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 12.200 7.700 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 8.600 4.300 12.200 10.100 ;
      RECT 3.400 11.500 9.600 12.500 ;
      RECT 8.600 4.300 9.600 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 8.600 16.300 12.200 19.700 ;
      RECT 0.800 18.700 12.200 19.700 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 8.600 28.300 9.600 29.300 ;
  END
END OR3FF

MACRO OR3GG
  CLASS CORE ;
  FOREIGN OR3GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 11.200 11.500 14.800 19.700 ;
      RECT 6.000 13.900 14.800 19.700 ;
      RECT 6.000 13.900 9.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 3.400 4.300 17.400 5.300 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 16.400 4.300 17.400 10.100 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 11.200 4.300 12.200 22.100 ;
      RECT 3.400 4.300 4.400 12.500 ;
      RECT 8.600 11.500 14.800 22.100 ;
      RECT 6.000 13.900 14.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 11.500 9.600 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OR3GG

MACRO OR3HH
  CLASS CORE ;
  FOREIGN OR3HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 20.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 17.300 ; # C|0.0@0
      RECT 0.800 16.300 4.400 17.300 ; # C|0.0@1
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 9.100 20.000 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 20.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 20.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 11.200 6.700 17.400 19.700 ;
      RECT 6.000 16.300 17.400 19.700 ;
      RECT 6.000 18.700 20.000 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 8.600 4.300 20.000 7.700 ;
      RECT 0.800 6.700 20.000 7.700 ;
      RECT 0.800 6.700 7.000 10.100 ;
      RECT 11.200 4.300 17.400 19.700 ;
      RECT 8.600 13.900 17.400 19.700 ;
      RECT 6.000 16.300 20.000 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 13.800 23.500 14.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END OR3HH

MACRO OR4EE
  CLASS CORE ;
  FOREIGN OR4EE 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 14.900 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 13.900 9.600 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 6.700 14.800 10.100 ; # Q|0.0@0
      RECT 13.800 13.900 14.800 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 10.100 ;
      RECT 3.400 11.500 14.800 12.500 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 12.200 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 9.600 12.500 ;
      RECT 13.800 4.300 14.800 12.500 ;
      RECT 0.800 6.700 14.800 12.500 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 11.200 16.300 14.800 19.700 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END OR4EE

MACRO OR4FF
  CLASS CORE ;
  FOREIGN OR4FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 12.500 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 6.700 14.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 0.800 18.700 12.200 19.700 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 9.600 0.500 ;
      RECT 0.800 4.300 4.400 7.700 ;
      RECT 8.600 4.300 9.600 7.700 ;
      RECT 13.800 4.300 14.800 7.700 ;
      RECT 0.800 6.700 14.800 7.700 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 0.800 11.500 12.200 12.500 ;
      RECT 0.800 16.300 1.800 19.700 ;
      RECT 11.200 16.300 14.800 19.700 ;
      RECT 0.800 18.700 14.800 19.700 ;
      RECT 13.800 16.300 14.800 22.100 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END OR4FF

MACRO OR4GG
  CLASS CORE ;
  FOREIGN OR4GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # D|0.0@0
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 11.200 6.700 12.200 19.700 ;
      RECT 11.200 13.900 14.800 19.700 ;
      RECT 8.600 16.300 14.800 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 0.800 4.300 17.400 5.300 ;
      RECT 3.400 4.300 12.200 7.700 ;
      RECT 16.400 4.300 17.400 10.100 ;
      RECT 3.400 4.300 4.400 10.100 ;
      RECT 11.200 4.300 12.200 19.700 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 11.500 7.000 14.900 ;
      RECT 6.000 13.900 14.800 14.900 ;
      RECT 8.600 13.900 14.800 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OR4GG

MACRO OR4HH
  CLASS CORE ;
  FOREIGN OR4HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 9.100 9.600 10.100 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 12.500 ; # C|0.0@0
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 19.700 ; # D|0.0@0
      RECT 0.800 18.700 14.800 19.700 ; # D|0.0@1
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 6.700 20.000 17.300 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 17.400 7.700 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 13.800 6.700 17.400 17.300 ;
      RECT 8.600 11.500 17.400 17.300 ;
      RECT 16.400 18.700 22.600 19.700 ;
      RECT 19.000 18.700 22.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 8.600 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 0.800 4.300 22.600 5.300 ;
      RECT 3.400 4.300 20.000 7.700 ;
      RECT 3.400 4.300 7.000 10.100 ;
      RECT 11.200 4.300 20.000 10.100 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 8.600 11.500 17.400 17.300 ;
      RECT 13.800 18.700 22.600 19.700 ;
      RECT 19.000 18.700 22.600 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 21.600 18.700 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END OR4HH

MACRO PDFF
  CLASS CORE ;
  FOREIGN PDFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END PDFF

MACRO PDGG
  CLASS CORE ;
  FOREIGN PDGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 0.800 9.100 1.800 10.100 ;
      RECT 3.400 11.500 4.400 14.900 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
  END
END PDGG

MACRO PUDD
  CLASS CORE ;
  FOREIGN PUDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 11.500 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 28.300 4.400 29.300 ;
  END
END PUDD

MACRO PUFF
  CLASS CORE ;
  FOREIGN PUFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 14.900 ; # Q|0.0@0
      RECT 0.800 13.900 4.400 14.900 ; # Q|0.0@1
      RECT 3.400 13.900 4.400 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 21.100 4.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 3.400 11.500 4.400 12.500 ;
      RECT 0.800 16.300 1.800 17.300 ;
      RECT 3.400 18.700 4.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END PUFF

MACRO PUGG
  CLASS CORE ;
  FOREIGN PUGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 7.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 9.100 4.400 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 14.900 ; # Q|0.0@0
      RECT 0.800 13.900 4.400 14.900 ; # Q|0.0@1
      RECT 3.400 13.900 4.400 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 7.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 7.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 3.400 11.500 4.400 12.500 ;
      RECT 0.800 16.300 4.400 17.300 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END PUGG

MACRO RSNDD
  CLASS CORE ;
  FOREIGN RSNDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # RN|0.0@0
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # SN|0.0@0
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 3.400 9.100 14.800 10.100 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 11.200 9.100 14.800 12.500 ;
      RECT 11.200 9.100 12.200 22.100 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 0.800 21.100 1.800 22.100 ;
      RECT 16.400 21.100 17.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 4.300 7.000 12.500 ;
      RECT 13.800 4.300 17.400 5.300 ;
      RECT 0.800 6.700 9.600 7.700 ;
      RECT 16.400 4.300 17.400 7.700 ;
      RECT 3.400 9.100 14.800 12.500 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 11.200 9.100 12.200 24.500 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 16.300 17.400 22.100 ;
      RECT 0.800 16.300 1.800 22.100 ;
      RECT 8.600 16.300 12.200 22.100 ;
      RECT 11.200 23.500 14.800 24.500 ;
      RECT 3.400 28.300 4.400 29.300 ;
  END
END RSNDD

MACRO SDCFF
  CLASS CORE ;
  FOREIGN SDCFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 67.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 13.900 33.000 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 13.900 12.200 14.900 ; # D|0.0@0
    END
  END D
  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 13.900 56.400 14.900 ; # CN|0.0@0
      RECT 6.000 16.300 7.000 19.700 ; # CN|0.0@1
      RECT 19.000 18.700 20.000 19.700 ; # CN|0.0@2
    END
  END CN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 11.500 20.000 14.900 ; # SI|0.0@0
    END
  END SI
  PIN T
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 22.100 ; # T|0.0@0
      RECT 58.000 9.100 59.000 10.100 ; # T|0.0@1
      RECT 55.400 16.300 59.000 17.300 ; # T|0.0@2
    END
  END T
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 65.800 6.700 66.800 7.700 ; # Q|0.0@0
      RECT 65.800 13.900 66.800 19.700 ; # Q|0.0@1
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 50.200 11.500 51.200 14.900 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 67.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 67.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 64.200 7.700 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 8.600 6.700 9.600 22.100 ;
      RECT 13.800 6.700 17.400 22.100 ;
      RECT 21.600 6.700 56.400 10.100 ;
      RECT 60.600 9.100 66.800 12.500 ;
      RECT 3.400 11.500 17.400 12.500 ;
      RECT 21.600 6.700 48.600 12.500 ;
      RECT 52.800 6.700 53.800 22.100 ;
      RECT 58.000 11.500 66.800 12.500 ;
      RECT 3.400 11.500 9.600 14.900 ;
      RECT 21.600 6.700 30.400 22.100 ;
      RECT 34.600 6.700 48.600 22.100 ;
      RECT 58.000 11.500 64.200 14.900 ;
      RECT 8.600 16.300 17.400 22.100 ;
      RECT 21.600 16.300 53.800 22.100 ;
      RECT 60.600 6.700 64.200 19.700 ;
      RECT 21.600 18.700 64.200 19.700 ;
      RECT 3.400 21.100 59.000 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 7.000 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 50.200 -0.500 51.200 0.500 ;
      RECT 55.400 -0.500 56.400 0.500 ;
      RECT 63.200 -0.500 64.200 0.500 ;
      RECT 0.800 4.300 56.400 5.300 ;
      RECT 63.200 4.300 66.800 14.900 ;
      RECT 0.800 4.300 1.800 7.700 ;
      RECT 6.000 6.700 66.800 7.700 ;
      RECT 6.000 4.300 17.400 12.500 ;
      RECT 21.600 4.300 40.800 12.500 ;
      RECT 45.000 4.300 56.400 10.100 ;
      RECT 60.600 6.700 66.800 14.900 ;
      RECT 0.800 11.500 40.800 12.500 ;
      RECT 45.000 4.300 48.600 12.500 ;
      RECT 52.800 11.500 66.800 12.500 ;
      RECT 3.400 11.500 9.600 14.900 ;
      RECT 13.800 4.300 17.400 24.500 ;
      RECT 21.600 4.300 30.400 24.500 ;
      RECT 34.600 4.300 40.800 24.500 ;
      RECT 47.600 4.300 48.600 24.500 ;
      RECT 52.800 4.300 53.800 24.500 ;
      RECT 58.000 11.500 66.800 14.900 ;
      RECT 3.400 11.500 4.400 24.500 ;
      RECT 8.600 16.300 17.400 24.500 ;
      RECT 21.600 16.300 53.800 24.500 ;
      RECT 60.600 6.700 64.200 19.700 ;
      RECT 21.600 18.700 66.800 19.700 ;
      RECT 3.400 21.100 59.000 22.100 ;
      RECT 65.800 18.700 66.800 22.100 ;
      RECT 0.800 23.500 56.400 24.500 ;
      RECT 63.200 23.500 64.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 14.800 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
      RECT 32.000 28.300 33.000 29.300 ;
      RECT 37.200 28.300 40.800 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 55.400 28.300 56.400 29.300 ;
      RECT 63.200 28.300 64.200 29.300 ;
  END
END SDCFF

MACRO SDFFFF
  CLASS CORE ;
  FOREIGN SDFFFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 52.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 11.500 14.800 14.900 ; # D|0.0@0
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 13.900 22.600 14.900 ; # SI|0.0@0
    END
  END SI
  PIN T
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 12.500 ; # T|0.0@0
    END
  END T
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 50.200 9.100 51.200 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 47.600 9.100 48.600 22.100 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 52.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 52.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 46.000 10.100 ;
      RECT 3.400 6.700 9.600 19.700 ;
      RECT 16.400 6.700 43.400 12.500 ;
      RECT 3.400 13.900 12.200 19.700 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 24.200 13.900 46.000 19.700 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 16.300 46.000 19.700 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 16.400 16.300 30.400 22.100 ;
      RECT 37.200 6.700 40.800 22.100 ;
      RECT 45.000 13.900 46.000 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 32.000 -0.500 35.600 0.500 ;
      RECT 42.400 -0.500 43.400 0.500 ;
      RECT 6.000 4.300 46.000 10.100 ;
      RECT 0.800 6.700 51.200 7.700 ;
      RECT 0.800 6.700 1.800 12.500 ;
      RECT 50.200 6.700 51.200 10.100 ;
      RECT 0.800 11.500 9.600 12.500 ;
      RECT 16.400 4.300 46.000 12.500 ;
      RECT 3.400 11.500 7.000 14.900 ;
      RECT 11.200 13.900 20.000 14.900 ;
      RECT 24.200 4.300 35.600 19.700 ;
      RECT 39.800 4.300 43.400 14.900 ;
      RECT 0.800 16.300 4.400 19.700 ;
      RECT 8.600 16.300 12.200 22.100 ;
      RECT 16.400 16.300 38.200 19.700 ;
      RECT 42.400 16.300 46.000 22.100 ;
      RECT 50.200 16.300 51.200 22.100 ;
      RECT 0.800 18.700 38.200 19.700 ;
      RECT 3.400 18.700 33.000 22.100 ;
      RECT 37.200 21.100 46.000 22.100 ;
      RECT 0.800 23.500 9.600 24.500 ;
      RECT 13.800 18.700 14.800 24.500 ;
      RECT 21.600 16.300 22.600 24.500 ;
      RECT 32.000 4.300 33.000 24.500 ;
      RECT 37.200 21.100 40.800 24.500 ;
      RECT 45.000 23.500 48.600 24.500 ;
      RECT 32.000 28.300 33.000 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
  END
END SDFFFF

MACRO SDPFF
  CLASS CORE ;
  FOREIGN SDPFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 75.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # CLK|0.0@0
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 12.500 ; # D|0.0@0
    END
  END D
  PIN PN
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 55.400 11.500 56.400 14.900 ; # PN|0.0@0
    END
  END PN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # SI|0.0@0
    END
  END SI
  PIN T
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 60.600 11.500 61.600 12.500 ; # T|0.0@0
    END
  END T
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 73.600 6.700 74.600 19.700 ; # Q|0.0@0
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 68.400 11.500 69.400 19.700 ; # QN|0.0@0
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 75.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 75.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 72.000 7.700 ;
      RECT 3.400 6.700 59.000 10.100 ;
      RECT 63.200 6.700 72.000 10.100 ;
      RECT 3.400 6.700 7.000 17.300 ;
      RECT 11.200 6.700 20.000 22.100 ;
      RECT 26.800 6.700 53.800 14.900 ;
      RECT 58.000 6.700 59.000 17.300 ;
      RECT 63.200 6.700 66.800 22.100 ;
      RECT 71.000 6.700 72.000 14.900 ;
      RECT 3.400 13.900 20.000 17.300 ;
      RECT 24.200 13.900 53.800 14.900 ;
      RECT 3.400 16.300 43.400 17.300 ;
      RECT 47.600 16.300 66.800 17.300 ;
      RECT 6.000 18.700 56.400 22.100 ;
      RECT 60.600 16.300 66.800 22.100 ;
      RECT 6.000 21.100 66.800 22.100 ;
      RECT 73.600 21.100 74.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 9.600 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 37.200 -0.500 38.200 0.500 ;
      RECT 42.400 -0.500 46.000 0.500 ;
      RECT 60.600 -0.500 61.600 0.500 ;
      RECT 65.800 -0.500 66.800 0.500 ;
      RECT 71.000 -0.500 72.000 0.500 ;
      RECT 0.800 4.300 74.600 5.300 ;
      RECT 3.400 4.300 69.400 7.700 ;
      RECT 73.600 4.300 74.600 10.100 ;
      RECT 0.800 9.100 46.000 10.100 ;
      RECT 50.200 4.300 69.400 10.100 ;
      RECT 0.800 9.100 7.000 12.500 ;
      RECT 11.200 4.300 20.000 24.500 ;
      RECT 26.800 11.500 53.800 12.500 ;
      RECT 58.000 4.300 59.000 12.500 ;
      RECT 63.200 4.300 66.800 24.500 ;
      RECT 71.000 11.500 72.000 14.900 ;
      RECT 3.400 13.900 51.200 14.900 ;
      RECT 60.600 13.900 66.800 19.700 ;
      RECT 3.400 4.300 4.400 17.300 ;
      RECT 8.600 13.900 43.400 24.500 ;
      RECT 47.600 11.500 51.200 19.700 ;
      RECT 55.400 16.300 69.400 19.700 ;
      RECT 73.600 16.300 74.600 22.100 ;
      RECT 8.600 18.700 69.400 19.700 ;
      RECT 3.400 21.100 48.600 22.100 ;
      RECT 52.800 18.700 56.400 22.100 ;
      RECT 63.200 16.300 69.400 22.100 ;
      RECT 0.800 23.500 43.400 24.500 ;
      RECT 47.600 11.500 48.600 24.500 ;
      RECT 71.000 23.500 72.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 12.200 29.300 ;
      RECT 34.600 28.300 40.800 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
      RECT 58.000 28.300 61.600 29.300 ;
      RECT 71.000 28.300 72.000 29.300 ;
  END
END SDPFF

MACRO THIGH
  CLASS CORE ;
  FOREIGN THIGH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN THIGH
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 13.900 4.400 17.300 ; # THIGH|0.0@0
    END
  END THIGH
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 18.700 4.400 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 3.400 16.300 4.400 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
  END
END THIGH

MACRO TLOW
  CLASS CORE ;
  FOREIGN TLOW 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 5.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN TLOW
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # TLOW|0.0@0
    END
  END TLOW
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 5.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 5.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 7.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 3.400 4.300 4.400 5.300 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 3.400 23.500 4.400 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
  END
END TLOW

MACRO TRIZDD
  FOREIGN TRIZDD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 13.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 13.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 13.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 10.100 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 8.600 6.700 9.600 19.700 ;
      RECT 3.400 13.900 9.600 17.300 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 3.400 4.300 9.600 7.700 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 3.400 4.300 7.000 10.100 ;
      RECT 11.200 6.700 12.200 12.500 ;
      RECT 0.800 11.500 4.400 12.500 ;
      RECT 8.600 11.500 12.200 12.500 ;
      RECT 3.400 13.900 9.600 17.300 ;
      RECT 3.400 16.300 12.200 17.300 ;
      RECT 3.400 4.300 4.400 22.100 ;
      RECT 8.600 11.500 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 8.600 23.500 9.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 8.600 28.300 9.600 29.300 ;
  END
END TRIZDD

MACRO TRIZFF
  CLASS CORE ;
  FOREIGN TRIZFF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 15.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 9.100 14.800 12.500 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 15.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 15.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 12.200 7.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 12.200 17.300 ;
      RECT 3.400 13.900 12.200 17.300 ;
      RECT 3.400 16.300 14.800 17.300 ;
      RECT 3.400 13.900 9.600 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 3.400 4.300 14.800 5.300 ;
      RECT 0.800 6.700 12.200 7.700 ;
      RECT 0.800 6.700 4.400 10.100 ;
      RECT 8.600 9.100 14.800 10.100 ;
      RECT 3.400 4.300 4.400 19.700 ;
      RECT 8.600 4.300 12.200 14.900 ;
      RECT 3.400 13.900 12.200 14.900 ;
      RECT 3.400 13.900 9.600 19.700 ;
      RECT 13.800 16.300 14.800 19.700 ;
      RECT 0.800 18.700 9.600 19.700 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
  END
END TRIZFF

MACRO TRIZGG
  CLASS CORE ;
  FOREIGN TRIZGG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 12.500 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 6.700 17.400 17.300 ; # Q|0.0@0
      RECT 13.800 18.700 14.800 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 14.800 7.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 14.800 10.100 ;
      RECT 8.600 6.700 12.200 22.100 ;
      RECT 8.600 13.900 14.800 17.300 ;
      RECT 3.400 18.700 12.200 19.700 ;
      RECT 8.600 21.100 17.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 7.000 0.500 ;
      RECT 3.400 4.300 17.400 10.100 ;
      RECT 3.400 4.300 4.400 22.100 ;
      RECT 8.600 4.300 12.200 24.500 ;
      RECT 0.800 13.900 14.800 14.900 ;
      RECT 3.400 13.900 14.800 22.100 ;
      RECT 3.400 18.700 17.400 22.100 ;
      RECT 6.000 18.700 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
  END
END TRIZGG

MACRO TRIZHH
  CLASS CORE ;
  FOREIGN TRIZHH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 23.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 11.500 22.600 14.900 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 9.100 1.800 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 11.200 11.500 12.200 14.900 ; # Q|0.0@0
      RECT 13.800 16.300 14.800 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 23.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 23.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 22.600 7.700 ;
      RECT 3.400 6.700 14.800 10.100 ;
      RECT 19.000 6.700 20.000 17.300 ;
      RECT 6.000 6.700 9.600 22.100 ;
      RECT 16.400 11.500 20.000 17.300 ;
      RECT 13.800 13.900 20.000 14.900 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 16.300 22.600 17.300 ;
      RECT 0.800 18.700 17.400 19.700 ;
      RECT 6.000 18.700 17.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 3.400 4.300 22.600 7.700 ;
      RECT 3.400 4.300 14.800 10.100 ;
      RECT 0.800 11.500 1.800 19.700 ;
      RECT 6.000 4.300 9.600 22.100 ;
      RECT 16.400 11.500 20.000 19.700 ;
      RECT 0.800 13.900 9.600 19.700 ;
      RECT 13.800 13.900 22.600 14.900 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 13.900 22.600 19.700 ;
      RECT 0.800 18.700 22.600 19.700 ;
      RECT 6.000 18.700 17.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 4.300 7.000 24.500 ;
      RECT 19.000 23.500 20.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 19.000 28.300 20.000 29.300 ;
  END
END TRIZHH

MACRO TRIZII
  CLASS CORE ;
  FOREIGN TRIZII 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 13.800 13.900 14.800 14.900 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 9.100 27.800 10.100 ; # Q|0.0@0
      RECT 21.600 9.100 22.600 14.900 ; # Q|0.0@1
      RECT 26.800 9.100 27.800 17.300 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 27.800 7.700 ;
      RECT 0.800 6.700 1.800 10.100 ;
      RECT 6.000 6.700 20.000 10.100 ;
      RECT 8.600 6.700 20.000 12.500 ;
      RECT 8.600 6.700 12.200 22.100 ;
      RECT 16.400 6.700 20.000 22.100 ;
      RECT 24.200 13.900 25.200 22.100 ;
      RECT 3.400 16.300 25.200 19.700 ;
      RECT 3.400 18.700 30.400 19.700 ;
      RECT 8.600 18.700 30.400 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 29.400 -0.500 30.400 0.500 ;
      RECT 0.800 4.300 25.200 7.700 ;
      RECT 0.800 6.700 27.800 7.700 ;
      RECT 0.800 4.300 1.800 10.100 ;
      RECT 6.000 4.300 20.000 12.500 ;
      RECT 26.800 6.700 27.800 10.100 ;
      RECT 24.200 11.500 25.200 22.100 ;
      RECT 8.600 4.300 12.200 22.100 ;
      RECT 16.400 4.300 20.000 22.100 ;
      RECT 3.400 16.300 27.800 22.100 ;
      RECT 3.400 18.700 30.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 16.300 7.000 24.500 ;
      RECT 13.800 16.300 14.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 13.800 28.300 14.800 29.300 ;
  END
END TRIZII

MACRO TRIZJJ
  CLASS CORE ;
  FOREIGN TRIZJJ 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 41.600 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 19.000 11.500 22.600 12.500 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 9.600 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 9.100 30.400 10.100 ; # Q|0.0@0
      RECT 37.200 9.100 38.200 17.300 ; # Q|0.0@1
      RECT 32.000 11.500 33.000 12.500 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 41.600 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 41.600 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 38.200 7.700 ;
      RECT 3.400 6.700 7.000 10.100 ;
      RECT 11.200 6.700 14.800 19.700 ;
      RECT 19.000 6.700 27.800 10.100 ;
      RECT 32.000 6.700 35.600 10.100 ;
      RECT 24.200 11.500 30.400 22.100 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 13.900 14.800 19.700 ;
      RECT 24.200 13.900 35.600 22.100 ;
      RECT 3.400 16.300 14.800 19.700 ;
      RECT 19.000 16.300 35.600 22.100 ;
      RECT 3.400 18.700 40.800 19.700 ;
      RECT 13.800 18.700 40.800 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 13.800 -0.500 14.800 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 39.800 -0.500 40.800 0.500 ;
      RECT 0.800 4.300 38.200 5.300 ;
      RECT 3.400 4.300 38.200 7.700 ;
      RECT 3.400 4.300 14.800 10.100 ;
      RECT 19.000 4.300 27.800 10.100 ;
      RECT 32.000 4.300 35.600 10.100 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 11.200 4.300 14.800 19.700 ;
      RECT 21.600 11.500 30.400 22.100 ;
      RECT 34.600 4.300 35.600 22.100 ;
      RECT 0.800 13.900 14.800 19.700 ;
      RECT 19.000 13.900 35.600 22.100 ;
      RECT 19.000 16.300 38.200 22.100 ;
      RECT 0.800 18.700 40.800 19.700 ;
      RECT 13.800 18.700 40.800 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 18.700 17.400 24.500 ;
      RECT 21.600 4.300 22.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
  END
END TRIZJJ

MACRO TRIZKK
  CLASS CORE ;
  FOREIGN TRIZKK 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 59.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 58.000 11.500 59.000 14.900 ; # E|0.0@0
    END
  END E
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 20.000 12.500 ; # A|0.0@0
    END
  END A
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 9.100 30.400 12.500 ; # Q|0.0@0
      RECT 42.400 9.100 43.400 17.300 ; # Q|0.0@1
      RECT 32.000 16.300 33.000 17.300 ; # Q|0.0@2
      RECT 37.200 16.300 38.200 17.300 ; # Q|0.0@3
      RECT 47.600 16.300 51.200 17.300 ; # Q|0.0@4
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 59.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 59.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 48.600 7.700 ;
      RECT 52.800 6.700 56.400 14.900 ;
      RECT 0.800 9.100 27.800 10.100 ;
      RECT 34.600 6.700 38.200 14.900 ;
      RECT 45.000 6.700 48.600 14.900 ;
      RECT 21.600 6.700 27.800 19.700 ;
      RECT 45.000 11.500 56.400 14.900 ;
      RECT 19.000 13.900 40.800 14.900 ;
      RECT 3.400 16.300 30.400 19.700 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 39.800 13.900 40.800 22.100 ;
      RECT 45.000 6.700 46.000 22.100 ;
      RECT 55.400 6.700 56.400 19.700 ;
      RECT 3.400 18.700 48.600 19.700 ;
      RECT 24.200 18.700 48.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 8.600 -0.500 9.600 0.500 ;
      RECT 16.400 -0.500 17.400 0.500 ;
      RECT 21.600 -0.500 22.600 0.500 ;
      RECT 50.200 -0.500 51.200 0.500 ;
      RECT 58.000 -0.500 59.000 0.500 ;
      RECT 0.800 4.300 59.000 5.300 ;
      RECT 3.400 4.300 48.600 7.700 ;
      RECT 52.800 4.300 56.400 10.100 ;
      RECT 0.800 9.100 30.400 10.100 ;
      RECT 34.600 4.300 38.200 14.900 ;
      RECT 42.400 4.300 48.600 10.100 ;
      RECT 6.000 4.300 7.000 19.700 ;
      RECT 13.800 4.300 14.800 19.700 ;
      RECT 21.600 4.300 27.800 19.700 ;
      RECT 45.000 11.500 53.800 14.900 ;
      RECT 3.400 13.900 40.800 14.900 ;
      RECT 45.000 13.900 59.000 14.900 ;
      RECT 3.400 13.900 30.400 19.700 ;
      RECT 34.600 4.300 35.600 22.100 ;
      RECT 39.800 13.900 40.800 22.100 ;
      RECT 45.000 4.300 46.000 22.100 ;
      RECT 50.200 11.500 51.200 17.300 ;
      RECT 55.400 13.900 56.400 22.100 ;
      RECT 3.400 18.700 48.600 19.700 ;
      RECT 24.200 18.700 48.600 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 23.500 7.000 24.500 ;
      RECT 11.200 23.500 12.200 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 24.200 4.300 25.200 24.500 ;
      RECT 52.800 23.500 53.800 24.500 ;
      RECT 58.000 23.500 59.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 11.200 28.300 12.200 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 52.800 28.300 53.800 29.300 ;
      RECT 58.000 28.300 59.000 29.300 ;
  END
END TRIZKK

MACRO XNOR2DD
  CLASS CORE ;
  FOREIGN XNOR2DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 13.900 17.400 17.300 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # Q|0.0@0
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 17.400 12.500 ;
      RECT 8.600 6.700 14.800 19.700 ;
      RECT 3.400 16.300 14.800 17.300 ;
      RECT 8.600 18.700 17.400 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 0.800 4.300 1.800 5.300 ;
      RECT 13.800 4.300 17.400 12.500 ;
      RECT 3.400 6.700 4.400 10.100 ;
      RECT 11.200 6.700 17.400 12.500 ;
      RECT 3.400 9.100 17.400 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 8.600 9.100 17.400 12.500 ;
      RECT 8.600 9.100 14.800 14.900 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 16.300 17.400 24.500 ;
      RECT 0.800 18.700 17.400 19.700 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 13.800 18.700 17.400 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
  END
END XNOR2DD

MACRO XNOR2FF
  CLASS CORE ;
  FOREIGN XNOR2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 11.500 17.400 17.300 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 17.400 7.700 ;
      RECT 3.400 6.700 14.800 10.100 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 8.600 6.700 14.800 22.100 ;
      RECT 3.400 16.300 14.800 22.100 ;
      RECT 3.400 18.700 17.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 13.800 -0.500 17.400 0.500 ;
      RECT 3.400 4.300 17.400 7.700 ;
      RECT 3.400 4.300 12.200 10.100 ;
      RECT 3.400 4.300 4.400 12.500 ;
      RECT 8.600 11.500 14.800 22.100 ;
      RECT 0.800 13.900 1.800 24.500 ;
      RECT 0.800 16.300 17.400 22.100 ;
      RECT 16.400 16.300 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END XNOR2FF

MACRO XNOR2GG
  CLASS CORE ;
  FOREIGN XNOR2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 13.900 27.800 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 9.600 12.500 ; # Q|0.0@0
      RECT 19.000 18.700 20.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 30.400 7.700 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 21.600 6.700 25.200 22.100 ;
      RECT 29.400 6.700 30.400 22.100 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 11.200 11.500 30.400 12.500 ;
      RECT 3.400 13.900 25.200 14.900 ;
      RECT 3.400 13.900 17.400 22.100 ;
      RECT 3.400 21.100 25.200 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 0.800 4.300 30.400 5.300 ;
      RECT 3.400 4.300 25.200 10.100 ;
      RECT 3.400 9.100 30.400 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 11.200 9.100 30.400 12.500 ;
      RECT 3.400 13.900 25.200 14.900 ;
      RECT 29.400 9.100 30.400 22.100 ;
      RECT 3.400 13.900 17.400 22.100 ;
      RECT 21.600 4.300 25.200 22.100 ;
      RECT 3.400 18.700 25.200 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 4.300 7.000 24.500 ;
      RECT 21.600 4.300 22.600 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END XNOR2GG

MACRO XNOR2HH
  CLASS CORE ;
  FOREIGN XNOR2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 36.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 11.500 33.000 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 20.000 12.500 ; # Q|0.0@0
      RECT 13.800 11.500 14.800 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 36.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 36.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 30.400 7.700 ;
      RECT 34.600 6.700 35.600 19.700 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 30.400 10.100 ;
      RECT 21.600 6.700 30.400 12.500 ;
      RECT 3.400 13.900 12.200 19.700 ;
      RECT 24.200 6.700 27.800 22.100 ;
      RECT 16.400 16.300 35.600 17.300 ;
      RECT 3.400 18.700 30.400 19.700 ;
      RECT 6.000 18.700 30.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 3.400 4.300 33.000 5.300 ;
      RECT 3.400 4.300 30.400 10.100 ;
      RECT 34.600 6.700 35.600 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 4.300 7.000 24.500 ;
      RECT 21.600 11.500 33.000 12.500 ;
      RECT 6.000 13.900 12.200 22.100 ;
      RECT 16.400 13.900 22.600 14.900 ;
      RECT 26.800 4.300 27.800 17.300 ;
      RECT 34.600 13.900 35.600 22.100 ;
      RECT 3.400 16.300 12.200 19.700 ;
      RECT 16.400 13.900 17.400 22.100 ;
      RECT 24.200 16.300 27.800 17.300 ;
      RECT 3.400 18.700 25.200 19.700 ;
      RECT 29.400 18.700 30.400 22.100 ;
      RECT 6.000 21.100 30.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 26.800 21.100 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 26.800 28.300 33.000 29.300 ;
  END
END XNOR2HH

MACRO XOR2DD
  CLASS CORE ;
  FOREIGN XOR2DD 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 13.900 17.400 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # Q|0.0@0
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 17.400 12.500 ;
      RECT 8.600 6.700 14.800 19.700 ;
      RECT 3.400 16.300 17.400 17.300 ;
      RECT 8.600 16.300 17.400 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 0.800 4.300 14.800 5.300 ;
      RECT 0.800 4.300 1.800 12.500 ;
      RECT 6.000 6.700 17.400 10.100 ;
      RECT 0.800 9.100 17.400 10.100 ;
      RECT 8.600 6.700 17.400 12.500 ;
      RECT 3.400 13.900 4.400 19.700 ;
      RECT 8.600 4.300 14.800 17.300 ;
      RECT 0.800 16.300 17.400 17.300 ;
      RECT 0.800 16.300 12.200 19.700 ;
      RECT 16.400 16.300 17.400 19.700 ;
      RECT 13.800 23.500 17.400 24.500 ;
      RECT 0.800 28.300 4.400 29.300 ;
  END
END XOR2DD

MACRO XOR2FF
  CLASS CORE ;
  FOREIGN XOR2FF 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 18.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 16.400 11.500 17.400 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 11.500 7.000 14.900 ; # Q|0.0@0
      RECT 6.000 18.700 7.000 19.700 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 18.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 18.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 0.800 6.700 17.400 10.100 ;
      RECT 3.400 6.700 4.400 19.700 ;
      RECT 8.600 6.700 14.800 19.700 ;
      RECT 3.400 16.300 17.400 17.300 ;
      RECT 8.600 16.300 17.400 19.700 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 11.200 -0.500 12.200 0.500 ;
      RECT 0.800 4.300 17.400 10.100 ;
      RECT 8.600 4.300 14.800 19.700 ;
      RECT 0.800 13.900 1.800 19.700 ;
      RECT 0.800 16.300 17.400 19.700 ;
      RECT 3.400 16.300 7.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 16.400 23.500 17.400 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 16.400 28.300 17.400 29.300 ;
  END
END XOR2FF

MACRO XOR2GG
  CLASS CORE ;
  FOREIGN XOR2GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 31.200 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 13.900 27.800 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 14.800 12.500 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 31.200 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 31.200 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 30.400 7.700 ;
      RECT 3.400 6.700 17.400 10.100 ;
      RECT 21.600 6.700 25.200 19.700 ;
      RECT 29.400 6.700 30.400 19.700 ;
      RECT 3.400 6.700 7.000 22.100 ;
      RECT 16.400 11.500 30.400 12.500 ;
      RECT 11.200 13.900 25.200 14.900 ;
      RECT 3.400 16.300 17.400 22.100 ;
      RECT 3.400 18.700 25.200 19.700 ;
      RECT 3.400 18.700 20.000 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 19.000 -0.500 20.000 0.500 ;
      RECT 0.800 4.300 30.400 5.300 ;
      RECT 3.400 4.300 30.400 7.700 ;
      RECT 3.400 4.300 17.400 10.100 ;
      RECT 21.600 4.300 30.400 10.100 ;
      RECT 0.800 11.500 7.000 12.500 ;
      RECT 19.000 11.500 27.800 12.500 ;
      RECT 3.400 13.900 25.200 14.900 ;
      RECT 29.400 13.900 30.400 19.700 ;
      RECT 3.400 13.900 17.400 22.100 ;
      RECT 21.600 4.300 25.200 19.700 ;
      RECT 3.400 18.700 25.200 19.700 ;
      RECT 3.400 18.700 20.000 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 6.000 4.300 7.000 24.500 ;
      RECT 21.600 23.500 22.600 24.500 ;
      RECT 26.800 23.500 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 26.800 28.300 27.800 29.300 ;
  END
END XOR2GG

MACRO XOR2HH
  CLASS CORE ;
  FOREIGN XOR2HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 36.400 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 11.500 1.800 14.900 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 32.000 11.500 33.000 14.900 ; # B|0.0@0
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 8.600 11.500 20.000 12.500 ; # Q|0.0@0
      RECT 13.800 11.500 14.800 17.300 ; # Q|0.0@1
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 36.400 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 36.400 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 30.400 7.700 ;
      RECT 34.600 6.700 35.600 22.100 ;
      RECT 3.400 6.700 4.400 22.100 ;
      RECT 8.600 6.700 30.400 10.100 ;
      RECT 21.600 6.700 30.400 12.500 ;
      RECT 3.400 13.900 12.200 22.100 ;
      RECT 24.200 6.700 30.400 22.100 ;
      RECT 16.400 16.300 35.600 19.700 ;
      RECT 3.400 18.700 35.600 19.700 ;
      RECT 3.400 18.700 30.400 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 4.400 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 32.000 -0.500 33.000 0.500 ;
      RECT 3.400 4.300 33.000 5.300 ;
      RECT 3.400 4.300 30.400 10.100 ;
      RECT 34.600 6.700 35.600 10.100 ;
      RECT 0.800 11.500 1.800 12.500 ;
      RECT 6.000 4.300 7.000 24.500 ;
      RECT 21.600 11.500 33.000 12.500 ;
      RECT 6.000 13.900 12.200 22.100 ;
      RECT 16.400 13.900 30.400 22.100 ;
      RECT 34.600 13.900 35.600 22.100 ;
      RECT 3.400 16.300 12.200 22.100 ;
      RECT 16.400 16.300 35.600 19.700 ;
      RECT 3.400 18.700 35.600 19.700 ;
      RECT 3.400 18.700 30.400 22.100 ;
      RECT 0.800 23.500 1.800 24.500 ;
      RECT 26.800 4.300 27.800 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 26.800 28.300 33.000 29.300 ;
  END
END XOR2HH

MACRO XOR3GG
  CLASS CORE ;
  FOREIGN XOR3GG 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 46.800 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 26.800 16.300 27.800 17.300 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 21.600 16.300 22.600 17.300 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 13.900 7.000 14.900 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.800 6.700 1.800 10.100 ; # Q|0.0@0
      RECT 0.800 9.100 4.400 10.100 ; # Q|0.0@1
      RECT 3.400 9.100 4.400 19.700 ; # Q|0.0@2
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 46.800 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 46.800 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 3.400 6.700 43.400 7.700 ;
      RECT 6.000 9.100 46.000 12.500 ;
      RECT 0.800 11.500 1.800 22.100 ;
      RECT 8.600 9.100 46.000 14.900 ;
      RECT 8.600 6.700 20.000 22.100 ;
      RECT 24.200 6.700 25.200 22.100 ;
      RECT 29.400 9.100 46.000 22.100 ;
      RECT 24.200 18.700 46.000 22.100 ;
      RECT 0.800 21.100 20.000 22.100 ;
    LAYER cont2 ;
      RECT 3.400 -0.500 4.400 0.500 ;
      RECT 21.600 -0.500 30.400 0.500 ;
      RECT 34.600 -0.500 35.600 0.500 ;
      RECT 42.400 -0.500 43.400 0.500 ;
      RECT 0.800 4.300 1.800 14.900 ;
      RECT 6.000 4.300 43.400 5.300 ;
      RECT 0.800 6.700 40.800 7.700 ;
      RECT 45.000 6.700 46.000 24.500 ;
      RECT 6.000 4.300 40.800 10.100 ;
      RECT 6.000 4.300 33.000 12.500 ;
      RECT 37.200 11.500 46.000 24.500 ;
      RECT 8.600 13.900 46.000 14.900 ;
      RECT 3.400 16.300 4.400 24.500 ;
      RECT 8.600 4.300 20.000 22.100 ;
      RECT 24.200 4.300 25.200 24.500 ;
      RECT 29.400 13.900 46.000 24.500 ;
      RECT 24.200 18.700 46.000 24.500 ;
      RECT 3.400 21.100 46.000 22.100 ;
      RECT 0.800 23.500 14.800 24.500 ;
      RECT 21.600 21.100 46.000 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 21.600 28.300 22.600 29.300 ;
      RECT 39.800 28.300 40.800 29.300 ;
  END
END XOR3GG

MACRO XOR3HH
  CLASS CORE ;
  FOREIGN XOR3HH 0.000 -4.800 ;
  ORIGIN 0.000 4.800 ;
  SIZE 52.000 BY 38.400 ;
  SYMMETRY X Y ;
  SITE CORE26 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 29.400 11.500 30.400 12.500 ; # A|0.0@0
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 24.200 11.500 25.200 12.500 ; # B|0.0@0
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 6.000 9.100 7.000 12.500 ; # C|0.0@0
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 3.400 6.700 4.400 19.700 ; # Q|0.0@0
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 23.600 52.000 29.200 ; # VDD|0.0@0
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    CAPACITANCE 0.00 ;
    PORT
    LAYER metal1 ;
      RECT 0.000 -0.400 52.000 5.200 ; # GND|0.0@0
    END
  END GND
  OBS
    LAYER metal1 ;
      RECT 8.600 6.700 51.200 10.100 ;
      RECT 0.800 11.500 1.800 22.100 ;
      RECT 8.600 6.700 22.600 17.300 ;
      RECT 26.800 6.700 27.800 22.100 ;
      RECT 32.000 6.700 51.200 17.300 ;
      RECT 8.600 13.900 51.200 17.300 ;
      RECT 13.800 6.700 22.600 22.100 ;
      RECT 26.800 13.900 46.000 22.100 ;
      RECT 0.800 21.100 22.600 22.100 ;
    LAYER cont2 ;
      RECT 0.800 -0.500 1.800 0.500 ;
      RECT 6.000 -0.500 7.000 0.500 ;
      RECT 24.200 -0.500 25.200 0.500 ;
      RECT 47.600 -0.500 48.600 0.500 ;
      RECT 3.400 4.300 4.400 7.700 ;
      RECT 8.600 4.300 51.200 7.700 ;
      RECT 8.600 4.300 48.600 10.100 ;
      RECT 0.800 11.500 1.800 14.900 ;
      RECT 6.000 11.500 22.600 12.500 ;
      RECT 26.800 4.300 27.800 17.300 ;
      RECT 39.800 11.500 51.200 17.300 ;
      RECT 8.600 13.900 30.400 17.300 ;
      RECT 37.200 13.900 51.200 17.300 ;
      RECT 3.400 16.300 4.400 24.500 ;
      RECT 8.600 16.300 51.200 17.300 ;
      RECT 13.800 4.300 22.600 22.100 ;
      RECT 29.400 16.300 46.000 24.500 ;
      RECT 3.400 21.100 22.600 22.100 ;
      RECT 26.800 21.100 46.000 24.500 ;
      RECT 0.800 23.500 17.400 24.500 ;
      RECT 24.200 23.500 48.600 24.500 ;
      RECT 0.800 28.300 1.800 29.300 ;
      RECT 6.000 28.300 7.000 29.300 ;
      RECT 24.200 28.300 25.200 29.300 ;
      RECT 47.600 28.300 48.600 29.300 ;
  END
END XOR3HH

MACRO PADCORNNE
FOREIGN PADCORNNE 0 0 ;
CLASS endcap topright ;
SITE necorner ;
SIZE 551.2 BY 551.2 ;
    OBS
        LAYER metal1 ; RECT 0 0 551.2 551.2 ;
        LAYER metal2 ; RECT 0 0 551.2 551.2 ;
        LAYER metal3 ; RECT 0 0 551.2 551.2 ;
    END
END PADCORNNE
MACRO PADCORNSE
FOREIGN PADCORNSE 0 0 ;
CLASS endcap bottomright ;
SITE secorner ;
SIZE 551.2 BY 551.2 ;
    OBS
        LAYER metal1 ; RECT 0 0 551.2 551.2 ;
        LAYER metal2 ; RECT 0 0 551.2 551.2 ;
        LAYER metal3 ; RECT 0 0 551.2 551.2 ;
    END
END PADCORNSE
MACRO PADCORNNW
FOREIGN PADCORNNW 0 0 ;
CLASS endcap topleft ;
SITE nwcorner ;
SIZE 551.2 BY 551.2 ;
    OBS
        LAYER metal1 ; RECT 0 0 551.2 551.2 ;
        LAYER metal2 ; RECT 0 0 551.2 551.2 ;
        LAYER metal3 ; RECT 0 0 551.2 551.2 ;
    END
END PADCORNNW
MACRO PADCORNSW
FOREIGN PADCORNSW 0 0 ;
CLASS endcap bottomleft ;
SITE swcorner ;
SIZE 551.2 BY 551.2 ;
   OBS
        LAYER metal1 ; RECT 0 0 551.2 551.2 ;
        LAYER metal2 ; RECT 0 0 551.2 551.2 ;
        LAYER metal3 ; RECT 0 0 551.2 551.2 ;
    END
END PADCORNSW
MACRO PADBGNDD
FOREIGN PADBGNDD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 5.2 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 5.2 551.2 ; RECT 0.0 0 4.2 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 5.2 551.2 ; RECT 0.0 0 4.2 2.3 ; 
      LAYER metal3 ; RECT 0 0 5.2 551.2 ;
      LAYER cont2 ; RECT 0 0 5.2 551.2 ;
      LAYER cont3 ; RECT 0 0 5.2 551.2 ;
   END
END PADBGNDD
MACRO PADBVDDD
FOREIGN PADBVDDD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 5.2 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 5.2 551.2 ; RECT 0.0 0 4.2 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 5.2 551.2 ; RECT 0.0 0 4.2 2.3 ; 
      LAYER metal3 ; RECT 0 0 5.2 551.2 ;
      LAYER cont2 ; RECT 0 0 5.2 551.2 ;
      LAYER cont3 ; RECT 0 0 5.2 551.2 ;
   END
END PADBVDDD
MACRO PADCINH0
FOREIGN PADCINH0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 43.7 2.3 ; RECT 47.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 43.7 2.3 ; RECT 47.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCINH0
MACRO PADCINH1
FOREIGN PADCINH1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCINH1
MACRO PADCINL0
FOREIGN PADCINL0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0370 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCINL0
MACRO PADCINL1
FOREIGN PADCINL1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCINL1
MACRO PADCIOH024
FOREIGN PADCIOH024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1060 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH024
MACRO PADCIOH024Q1
FOREIGN PADCIOH024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1060 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH024Q1
MACRO PADCIOH04
FOREIGN PADCIOH04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2230 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3800 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH04
MACRO PADCIOH08
FOREIGN PADCIOH08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0910 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH08
MACRO PADCIOH08F
FOREIGN PADCIOH08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5830 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2510 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 38.5 2.3 ; RECT 42.1 0 43.7 2.3 ;RECT 47.3 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH08F
MACRO PADCIOH124
FOREIGN PADCIOH124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1020 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1530 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH124
MACRO PADCIOH124Q1
FOREIGN PADCIOH124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1080 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH124Q1
MACRO PADCIOH14
FOREIGN PADCIOH14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2200 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3830 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH14
MACRO PADCIOH18
FOREIGN PADCIOH18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0630 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0930 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH18
MACRO PADCIOH18F
FOREIGN PADCIOH18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5850 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 44.7 0 46.3 1.3 ;
         LAYER metal2 ; RECT 44.7 0 46.3 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0300 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 43.7 2.3 ;RECT 47.3 0 48.9 2.3 ;RECT 52.5 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOH18F
MACRO PADCIOL024
FOREIGN PADCIOL024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1070 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1380 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0360 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL024
MACRO PADCIOL024Q1
FOREIGN PADCIOL024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0730 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0930 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0360 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL024Q1
MACRO PADCIOL04
FOREIGN PADCIOL04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2250 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0360 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL04
MACRO PADCIOL08
FOREIGN PADCIOL08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0360 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL08
MACRO PADCIOL08F
FOREIGN PADCIOL08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4280 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0360 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1540 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 33.3 2.3 ;RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL08F
MACRO PADCIOL124
FOREIGN PADCIOL124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1040 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1400 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL124
MACRO PADCIOL124Q1
FOREIGN PADCIOL124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0700 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0950 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL124Q1
MACRO PADCIOL14
FOREIGN PADCIOL14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL14
MACRO PADCIOL18
FOREIGN PADCIOL18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0800 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL18
MACRO PADCIOL18F
FOREIGN PADCIOL18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4250 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 39.5 0 41.1 1.3 ;
         LAYER metal2 ; RECT 39.5 0 41.1 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 100.9 1.3 ;
         LAYER metal2 ; RECT 96.7 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 10.9 0 38.5 2.3 ;RECT 42.1 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADCIOL18F
MACRO PADGNDD
FOREIGN PADGNDD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADGNDD
MACRO PADGNDIO
FOREIGN PADGNDIO 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADGNDIO
MACRO PADGNDIOD
FOREIGN PADGNDIOD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADGNDIOD
MACRO PADGNDIOL
FOREIGN PADGNDIOL 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN GND
      DIRECTION input ;
      CAPACITANCE 0.0000 ;
      USE ground ;
      PORT
         LAYER metal1 ; RECT 8.3 0 100.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 100.9 1.3 ;
      END
   END GND
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADGNDIOL
MACRO PADGNDL
FOREIGN PADGNDL 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN GND
      DIRECTION input ;
      CAPACITANCE 0.0000 ;
      USE ground ;
      PORT
         LAYER metal1 ; RECT 8.3 0 100.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 100.9 1.3 ;
      END
   END GND
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADGNDL
MACRO PADOUT16
FOREIGN PADOUT16 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0610 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0820 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADOUT16
MACRO PADOUT24
FOREIGN PADOUT24 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1000 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADOUT24
MACRO PADOUT4
FOREIGN PADOUT4 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2180 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3700 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADOUT4
MACRO PADOUT8
FOREIGN PADOUT8 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0610 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0810 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADOUT8
MACRO PADOUT8F
FOREIGN PADOUT8F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4210 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5730 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 46.3 2.3 ;RECT 49.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADOUT8F
MACRO PADSINH0
FOREIGN PADSINH0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.1790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 56.7 2.3 ; RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 56.7 2.3 ; RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSINH0
MACRO PADSINH1
FOREIGN PADSINH1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 56.7 2.3 ; RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 56.7 2.3 ; RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSINH1
MACRO PADSINL0
FOREIGN PADSINL0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 64.5 2.3 ; RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 64.5 2.3 ; RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSINL0
MACRO PADSINL1
FOREIGN PADSINL1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0250 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 64.5 2.3 ; RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 64.5 2.3 ; RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSINL1
MACRO PADSIOH024
FOREIGN PADSIOH024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1020 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.1790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH024
MACRO PADSIOH024Q1
FOREIGN PADSIOH024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0960 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.1790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH024Q1
MACRO PADSIOH04
FOREIGN PADSIOH04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2190 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.1790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH04
MACRO PADSIOH08
FOREIGN PADSIOH08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0630 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0820 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.1790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH08
MACRO PADSIOH08F
FOREIGN PADSIOH08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5730 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0000 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH08F
MACRO PADSIOH124
FOREIGN PADSIOH124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1010 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1410 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH124
MACRO PADSIOH124Q1
FOREIGN PADSIOH124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0960 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH124Q1
MACRO PADSIOH14
FOREIGN PADSIOH14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2190 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH14
MACRO PADSIOH18
FOREIGN PADSIOH18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0630 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0820 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH18
MACRO PADSIOH18F
FOREIGN PADSIOH18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5730 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0260 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2430 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 56.7 2.3 ;RECT 60.3 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOH18F
MACRO PADSIOL024
FOREIGN PADSIOL024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1020 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1450 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL024
MACRO PADSIOL024Q1
FOREIGN PADSIOL024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1000 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL024Q1
MACRO PADSIOL04
FOREIGN PADSIOL04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2200 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3740 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL04
MACRO PADSIOL08
FOREIGN PADSIOL08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0630 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0850 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL08
MACRO PADSIOL08F
FOREIGN PADSIOL08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0650 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL08F
MACRO PADSIOL124
FOREIGN PADSIOL124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1010 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1440 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0240 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL124
MACRO PADSIOL124Q1
FOREIGN PADSIOL124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0990 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0240 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL124Q1
MACRO PADSIOL14
FOREIGN PADSIOL14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2190 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3740 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0240 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL14
MACRO PADSIOL18
FOREIGN PADSIOL18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0620 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0840 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0250 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL18
MACRO PADSIOL18F
FOREIGN PADSIOL18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4210 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 52.5 0 54.1 1.3 ;
         LAYER metal2 ; RECT 52.5 0 54.1 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5760 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 34.3 0 35.9 1.3 ;
         LAYER metal2 ; RECT 34.3 0 35.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0240 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 65.5 0 67.1 1.3 ;
         LAYER metal2 ; RECT 65.5 0 67.1 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 98.3 1.3 ;
         LAYER metal2 ; RECT 94.1 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 33.3 2.3 ; RECT 36.9 0 51.5 2.3 ;RECT 55.1 0 64.5 2.3 ;RECT 68.1 0 93.1 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADSIOL18F
MACRO PADTCLH
FOREIGN PADTCLH 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.6290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 98.3 2.3 ; RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 98.3 2.3 ; RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTCLH
MACRO PADTCLH0
FOREIGN PADTCLH0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0900 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 60.3 0 61.9 1.3 ;
         LAYER metal2 ; RECT 60.3 0 61.9 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.6290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 59.3 2.3 ; RECT 62.9 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 59.3 2.3 ; RECT 62.9 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTCLH0
MACRO PADTINH0
FOREIGN PADTINH0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTINH0
MACRO PADTINH1
FOREIGN PADTINH1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2520 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTINH1
MACRO PADTINL0
FOREIGN PADTINL0 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTINL0
MACRO PADTINL1
FOREIGN PADTINL1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTINL1
MACRO PADTIOH016
FOREIGN PADTIOH016 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0620 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0840 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH016
MACRO PADTIOH024
FOREIGN PADTIOH024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1010 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1420 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH024
MACRO PADTIOH024Q1
FOREIGN PADTIOH024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0970 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH024Q1
MACRO PADTIOH04
FOREIGN PADTIOH04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2190 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3720 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH04
MACRO PADTIOH08
FOREIGN PADTIOH08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0620 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0830 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2490 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH08
MACRO PADTIOH08F
FOREIGN PADTIOH08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4220 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5750 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 5.7 0 7.3 1.3 ;
         LAYER metal2 ; RECT 5.7 0 7.3 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2500 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 94.1 0 100.9 1.3 ;
         LAYER metal2 ; RECT 94.1 0 100.9 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 4.7 2.3 ; RECT 8.3 0 15.1 2.3 ;RECT 18.7 0 46.3 2.3 ;RECT 49.9 0 93.1 2.3 ;RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH08F
MACRO PADTIOH124
FOREIGN PADTIOH124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1010 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1440 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2520 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH124
MACRO PADTIOH124Q1
FOREIGN PADTIOH124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0990 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2520 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH124Q1
MACRO PADTIOH14
FOREIGN PADTIOH14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2190 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3730 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2520 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH14
MACRO PADTIOH18
FOREIGN PADTIOH18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0620 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0840 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2530 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH18
MACRO PADTIOH18F
FOREIGN PADTIOH18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4210 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5760 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 8.3 0 9.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 9.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.2520 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 99.3 0 106.1 1.3 ;
         LAYER metal2 ; RECT 99.3 0 106.1 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 7.3 2.3 ;RECT 10.9 0 48.9 2.3 ;RECT 52.5 0 98.3 2.3 ;RECT 107.1 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOH18F
MACRO PADTIOL024
FOREIGN PADTIOL024 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1030 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1370 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 42.1 0 43.7 1.3 ;
         LAYER metal2 ; RECT 42.1 0 43.7 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL024
MACRO PADTIOL024Q1
FOREIGN PADTIOL024Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0920 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 42.1 0 43.7 1.3 ;
         LAYER metal2 ; RECT 42.1 0 43.7 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL024Q1
MACRO PADTIOL04
FOREIGN PADTIOL04 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2210 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 42.1 0 43.7 1.3 ;
         LAYER metal2 ; RECT 42.1 0 43.7 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL04
MACRO PADTIOL08
FOREIGN PADTIOL08 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0640 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0780 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 42.1 0 43.7 1.3 ;
         LAYER metal2 ; RECT 42.1 0 43.7 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL08
MACRO PADTIOL08F
FOREIGN PADTIOL08F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4240 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 49.9 0 51.5 1.3 ;
         LAYER metal2 ; RECT 49.9 0 51.5 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5690 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 42.1 0 43.7 1.3 ;
         LAYER metal2 ; RECT 42.1 0 43.7 1.3 ;
      END
   END O
   PIN IEN
      DIRECTION input ;
      CAPACITANCE 0.0680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 16.1 0 17.7 1.3 ;
         LAYER metal2 ; RECT 16.1 0 17.7 1.3 ;
      END
   END IEN
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1670 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 91.5 0 98.3 1.3 ;
         LAYER metal2 ; RECT 91.5 0 98.3 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 15.1 2.3 ; RECT 18.7 0 41.1 2.3 ;RECT 44.7 0 48.9 2.3 ;RECT 52.5 0 90.5 2.3 ;RECT 99.3 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL08F
MACRO PADTIOL124
FOREIGN PADTIOL124 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.1050 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.1380 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL124
MACRO PADTIOL124Q1
FOREIGN PADTIOL124Q1 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0710 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0930 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL124Q1
MACRO PADTIOL14
FOREIGN PADTIOL14 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.2230 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.3680 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL14
MACRO PADTIOL18
FOREIGN PADTIOL18 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.0660 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.0790 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL18
MACRO PADTIOL18F
FOREIGN PADTIOL18F 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN OEN
      DIRECTION input ;
      CAPACITANCE 0.4250 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 57.7 0 59.3 1.3 ;
         LAYER metal2 ; RECT 57.7 0 59.3 1.3 ;
      END
   END OEN
   PIN O
      DIRECTION input ;
      CAPACITANCE 0.5700 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 47.3 0 48.9 1.3 ;
         LAYER metal2 ; RECT 47.3 0 48.9 1.3 ;
      END
   END O
   PIN IE
      DIRECTION input ;
      CAPACITANCE 0.0290 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 3.1 0 4.7 1.3 ;
         LAYER metal2 ; RECT 3.1 0 4.7 1.3 ;
      END
   END IE
   PIN I
      DIRECTION output ;
      CAPACITANCE 0.1770 ;
      USE signal ;
      PORT
         LAYER metal1 ; RECT 96.7 0 103.5 1.3 ;
         LAYER metal2 ; RECT 96.7 0 103.5 1.3 ;
      END
   END I
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 2.1 2.3 ; RECT 5.7 0 46.3 2.3 ;RECT 49.9 0 56.7 2.3 ;RECT 60.3 0 95.7 2.3 ;RECT 104.5 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADTIOL18F
MACRO PADVDDD
FOREIGN PADVDDD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADVDDD
MACRO PADVDDIO
FOREIGN PADVDDIO 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADVDDIO
MACRO PADVDDIOD
FOREIGN PADVDDIOD 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 118.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADVDDIOD
MACRO PADVDDIOL
FOREIGN PADVDDIOL 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN VDD
      DIRECTION input ;
      CAPACITANCE 0.0000 ;
      USE power ;
      PORT
         LAYER metal1 ; RECT 8.3 0 100.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 100.9 1.3 ;
      END
   END VDD
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADVDDIOL
MACRO PADVDDL
FOREIGN PADVDDL 0 0 ;
CLASS pad ;
SITE target ;
SYMMETRY r90 ;
SIZE 119.6 by 551.2 ;
   PIN SIGNAME
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END SIGNAME
   PIN GEN
      DIRECTION inout ;
      CAPACITANCE 0 ;
      USE signal ;
      PORT
         # No port geometry defined ( unrouted signal )
      END
   END GEN
   PIN VDD
      DIRECTION input ;
      CAPACITANCE 0.0000 ;
      USE power ;
      PORT
         LAYER metal1 ; RECT 8.3 0 100.9 1.3 ;
         LAYER metal2 ; RECT 8.3 0 100.9 1.3 ;
      END
   END VDD
   OBS
      LAYER metal1 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal2 ; RECT 0 2.3 119.6 551.2 ; RECT 0.0 0 7.3 2.3 ; RECT 101.9 0 119.6 2.3 ; 
      LAYER metal3 ; RECT 0 0 119.6 551.2 ;
      LAYER cont2 ; RECT 0 0 119.6 551.2 ;
      LAYER cont3 ; RECT 0 0 119.6 551.2 ;
   END
END PADVDDL
MACRO ZZPADSPC
FOREIGN ZZPADSPC 0 0 ;
SYMMETRY r90 ;
CLASS pad ;
SITE target ;
SIZE 5.2 BY 551.2 ;
    OBS
        LAYER metal1 ; RECT 0 0 5.2 551.2 ;
        LAYER metal2 ; RECT 0 0 5.2 551.2 ;
        LAYER metal3 ; RECT 0 0 5.2 551.2 ;
    END
END ZZPADSPC

END LIBRARY
# /mnts/hpdtctm/cbs1/D3.1X/700/bin/gridit:
# 	 set-b.ada 1.6 93/05/05 15:24:33
# 	 attr_utils-s.ada 1.6 91/10/25 16:05:35 
# 	 attr_utils-b.ada 1.11 91/10/25 16:06:40 
# 	 coral_util-s.ada 1.19 92/09/02 11:27:39 
# 	 coral_util-b.ada 11.9 93/06/28 15:47:02 
# 	 datetime-b.ada 1.6 93/05/05 15:24:23
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 coral 12.2 92/10/12 10:58:44
# 	 dftogds-b.ada 1.10 93/05/24 15:37:06 
# 	 dstring-s.ada 11.2 93/05/05 15:24:29
# 	 set-b.ada 1.6 93/05/05 15:24:33
# 	 dstring-b.ada 11.2 93/05/05 15:24:27 
# 	 gdstodf-b.ada 1.7 93/05/05 15:27:04 
# 	 gridit-d.ada 1.11 93/05/24 15:37:10 
# 	 grid-b.ada 1.6 93/05/05 15:27:08 
# /mnts/hpdtctm/cbs1/D3.1X/700/bin/c3lefgen:
# 	 set-b.ada 1.6 93/05/05 15:24:33
# 	 attr_utils-s.ada 1.6 91/10/25 16:05:35 
# 	 attr_utils-b.ada 1.11 91/10/25 16:06:40 
# 	 bdltodf-b.ada 12.5 92/12/15 17:32:09 
# 	 bb_trees-b.ada 1.5 93/05/05 15:22:02
# 	 string_hash-b.ada 1.6 93/05/05 15:27:29 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 string_hash-s.ada 1.6 93/05/05 15:27:30 
# 	 bb_trees-b.ada 1.5 93/05/05 15:22:02
# 	 coral_hash-b.ada 1.4 93/05/05 15:27:22 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 coral_hash-s.ada 1.5 93/05/05 15:27:23 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 c3lefgen-d.ada 1.38 93/06/28 15:46:53 
# 	 coral_util-s.ada 1.19 92/09/02 11:27:39 
# 	 coral_util-b.ada 11.9 93/06/28 15:47:02 
# 	 data_file-b.ada 1.7 93/05/24 15:36:52 
# 	 datetime-b.ada 1.6 93/05/05 15:24:23
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 coral 12.2 92/10/12 10:58:44
# 	 dftobm-b.ada 1.37 93/06/28 15:47:06 
# 	 dftogds-b.ada 1.10 93/05/24 15:37:06 
# 	 dftolef-b.ada 12.18 93/06/28 15:47:08 
# 	 dstring-s.ada 11.2 93/05/05 15:24:29
# 	 set-b.ada 1.6 93/05/05 15:24:33
# 	 dstring-b.ada 11.2 93/05/05 15:24:27 
# 	 gdstodf-b.ada 1.7 93/05/05 15:27:04 
# 	 get_data-b.ada 1.10 93/05/24 15:36:54 
# 	 string_hash-b.ada 1.6 93/05/05 15:27:29 
# 	 map-s.ada 1.6 93/05/05 15:27:26 
# 	 string_hash-s.ada 1.6 93/05/05 15:27:30 
# 	 map-b.ada 1.7 93/05/05 15:27:25 
# 	 prim-b.ada 1.36 93/05/05 15:27:32 
# 	TAG: RELEASE_B_03_00                        
# 	 DFACCESS07  B.03.00 DF ACCESS ROUTINES                       17May93 
# 	Copyright Hewlett-Packard Co. 1992,1993                                
# 	 MP:	 KDFACCESS  0.09  17May93 15:41:16   

